magic
tech sky130A
timestamp 1697426997
<< nwell >>
rect -68 2495 1201 2496
rect -90 2491 1257 2495
rect -116 1716 1257 2491
<< nmos >>
rect 81 1301 131 1602
rect 181 1301 231 1602
rect 281 1301 351 1602
rect 401 1301 451 1602
rect 501 1301 551 1602
rect 601 1301 651 1602
rect 701 1301 751 1602
rect 801 1301 861 1602
rect 911 1301 961 1602
rect 1011 1301 1061 1602
rect 15 450 65 1050
rect 115 450 165 1050
rect 215 450 265 1050
rect 401 451 451 1051
rect 501 451 551 1051
rect 601 451 651 1051
rect 701 451 751 1051
rect 880 451 930 1051
rect 980 451 1030 1051
rect 1080 451 1130 1051
rect 15 -350 65 250
rect 115 -350 165 250
rect 215 -350 265 250
rect 401 -349 451 251
rect 501 -349 551 251
rect 601 -349 651 251
rect 701 -349 751 251
rect 880 -349 930 251
rect 980 -349 1030 251
rect 1080 -349 1130 251
<< pmos >>
rect 15 1806 65 2406
rect 115 1806 165 2406
rect 215 1806 265 2406
rect 401 1807 451 2407
rect 501 1807 551 2407
rect 601 1807 651 2407
rect 701 1807 751 2407
rect 880 1807 930 2407
rect 980 1807 1030 2407
rect 1080 1807 1130 2407
<< ndiff >>
rect 245 1602 267 1603
rect 465 1602 487 1603
rect 565 1602 587 1603
rect 31 1598 81 1602
rect 31 1316 46 1598
rect 66 1316 81 1598
rect 31 1301 81 1316
rect 131 1597 181 1602
rect 131 1316 146 1597
rect 166 1316 181 1597
rect 131 1301 181 1316
rect 231 1598 281 1602
rect 231 1316 246 1598
rect 266 1316 281 1598
rect 231 1301 281 1316
rect 351 1597 401 1602
rect 351 1316 366 1597
rect 386 1316 401 1597
rect 351 1301 401 1316
rect 451 1598 501 1602
rect 451 1316 466 1598
rect 486 1316 501 1598
rect 451 1301 501 1316
rect 551 1598 601 1602
rect 551 1316 566 1598
rect 586 1316 601 1598
rect 551 1301 601 1316
rect 651 1597 701 1602
rect 651 1316 666 1597
rect 686 1316 701 1597
rect 651 1301 701 1316
rect 751 1597 801 1602
rect 751 1316 766 1597
rect 786 1316 801 1597
rect 751 1301 801 1316
rect 861 1597 911 1602
rect 861 1316 876 1597
rect 896 1316 911 1597
rect 861 1301 911 1316
rect 961 1597 1011 1602
rect 961 1316 976 1597
rect 996 1316 1011 1597
rect 961 1301 1011 1316
rect 1061 1597 1109 1602
rect 1061 1316 1076 1597
rect 1096 1316 1109 1597
rect 1061 1301 1109 1316
rect -35 1035 15 1050
rect -35 470 -15 1035
rect 2 470 15 1035
rect -35 450 15 470
rect 65 1040 115 1050
rect 65 465 80 1040
rect 100 465 115 1040
rect 65 450 115 465
rect 165 1040 215 1050
rect 165 465 180 1040
rect 200 465 215 1040
rect 165 450 215 465
rect 265 1040 315 1050
rect 265 465 280 1040
rect 300 465 315 1040
rect 265 450 315 465
rect 351 1041 401 1051
rect 351 466 366 1041
rect 386 466 401 1041
rect 351 451 401 466
rect 451 1041 501 1051
rect 451 466 466 1041
rect 486 466 501 1041
rect 451 451 501 466
rect 551 1041 601 1051
rect 551 466 566 1041
rect 586 466 601 1041
rect 551 451 601 466
rect 651 1041 701 1051
rect 651 466 666 1041
rect 686 466 701 1041
rect 651 451 701 466
rect 751 1041 799 1051
rect 751 466 766 1041
rect 786 466 799 1041
rect 751 451 799 466
rect 830 1036 880 1051
rect 830 461 845 1036
rect 865 461 880 1036
rect 830 451 880 461
rect 930 1036 980 1051
rect 930 461 945 1036
rect 965 461 980 1036
rect 930 451 980 461
rect 1030 1036 1080 1051
rect 1030 461 1045 1036
rect 1065 461 1080 1036
rect 1030 451 1080 461
rect 1130 1036 1180 1051
rect 1130 461 1143 1036
rect 1163 461 1180 1036
rect 1130 451 1180 461
rect -35 240 15 250
rect -35 -335 -20 240
rect 0 -335 15 240
rect -35 -350 15 -335
rect 65 240 115 250
rect 65 -335 80 240
rect 100 -335 115 240
rect 65 -350 115 -335
rect 165 240 215 250
rect 165 -335 180 240
rect 200 -335 215 240
rect 165 -350 215 -335
rect 265 240 315 250
rect 265 -335 280 240
rect 300 -335 315 240
rect 265 -350 315 -335
rect 351 241 401 251
rect 351 -334 366 241
rect 386 -334 401 241
rect 351 -349 401 -334
rect 451 241 501 251
rect 451 -334 466 241
rect 486 -334 501 241
rect 451 -349 501 -334
rect 551 241 601 251
rect 551 -334 566 241
rect 586 -334 601 241
rect 551 -349 601 -334
rect 651 241 701 251
rect 651 -334 666 241
rect 686 -334 701 241
rect 651 -349 701 -334
rect 751 241 799 251
rect 751 -334 766 241
rect 786 -334 799 241
rect 751 -349 799 -334
rect 830 236 880 251
rect 830 -339 845 236
rect 865 -339 880 236
rect 830 -349 880 -339
rect 930 236 980 251
rect 930 -339 945 236
rect 965 -339 980 236
rect 930 -349 980 -339
rect 1030 236 1080 251
rect 1030 -339 1045 236
rect 1065 -339 1080 236
rect 1030 -349 1080 -339
rect 1130 236 1180 251
rect 1130 -339 1145 236
rect 1165 -339 1180 236
rect 1130 -349 1180 -339
<< pdiff >>
rect -35 2396 15 2406
rect -35 1821 -20 2396
rect 0 1821 15 2396
rect -35 1806 15 1821
rect 65 2396 115 2406
rect 65 1821 80 2396
rect 100 1821 115 2396
rect 65 1806 115 1821
rect 165 2396 215 2406
rect 165 1821 180 2396
rect 200 1821 215 2396
rect 165 1806 215 1821
rect 265 2396 315 2406
rect 265 1821 280 2396
rect 300 1821 315 2396
rect 265 1806 315 1821
rect 351 2397 401 2407
rect 351 1822 366 2397
rect 386 1822 401 2397
rect 351 1807 401 1822
rect 451 2397 501 2407
rect 451 1822 466 2397
rect 486 1822 501 2397
rect 451 1807 501 1822
rect 551 2397 601 2407
rect 551 1822 566 2397
rect 586 1822 601 2397
rect 551 1807 601 1822
rect 651 2397 701 2407
rect 651 1822 666 2397
rect 686 1822 701 2397
rect 651 1807 701 1822
rect 751 2397 799 2407
rect 751 1822 766 2397
rect 786 1822 799 2397
rect 751 1807 799 1822
rect 830 2392 880 2407
rect 830 1817 845 2392
rect 865 1817 880 2392
rect 830 1807 880 1817
rect 930 2392 980 2407
rect 930 1817 945 2392
rect 965 1817 980 2392
rect 930 1807 980 1817
rect 1030 2392 1080 2407
rect 1030 1817 1045 2392
rect 1065 1817 1080 2392
rect 1030 1807 1080 1817
rect 1130 2392 1180 2407
rect 1130 1817 1145 2392
rect 1165 1817 1180 2392
rect 1130 1807 1180 1817
<< ndiffc >>
rect 46 1316 66 1598
rect 146 1316 166 1597
rect 246 1316 266 1598
rect 366 1316 386 1597
rect 466 1316 486 1598
rect 566 1316 586 1598
rect 666 1316 686 1597
rect 766 1316 786 1597
rect 876 1316 896 1597
rect 976 1316 996 1597
rect 1076 1316 1096 1597
rect -15 470 2 1035
rect 80 465 100 1040
rect 180 465 200 1040
rect 280 465 300 1040
rect 366 466 386 1041
rect 466 466 486 1041
rect 566 466 586 1041
rect 666 466 686 1041
rect 766 466 786 1041
rect 845 461 865 1036
rect 945 461 965 1036
rect 1045 461 1065 1036
rect 1143 461 1163 1036
rect -20 -335 0 240
rect 80 -335 100 240
rect 180 -335 200 240
rect 280 -335 300 240
rect 366 -334 386 241
rect 466 -334 486 241
rect 566 -334 586 241
rect 666 -334 686 241
rect 766 -334 786 241
rect 845 -339 865 236
rect 945 -339 965 236
rect 1045 -339 1065 236
rect 1145 -339 1165 236
<< pdiffc >>
rect -20 1821 0 2396
rect 80 1821 100 2396
rect 180 1821 200 2396
rect 280 1821 300 2396
rect 366 1822 386 2397
rect 466 1822 486 2397
rect 566 1822 586 2397
rect 666 1822 686 2397
rect 766 1822 786 2397
rect 845 1817 865 2392
rect 945 1817 965 2392
rect 1045 1817 1065 2392
rect 1145 1817 1165 2392
<< psubdiff >>
rect 401 1191 446 1206
rect 401 1116 414 1191
rect 431 1116 446 1191
rect 401 1099 446 1116
rect 751 1191 796 1206
rect 751 1116 764 1191
rect 781 1116 796 1191
rect 751 1099 796 1116
<< nsubdiff >>
rect -85 2392 -35 2406
rect -85 1822 -70 2392
rect -44 1822 -35 2392
rect -85 1806 -35 1822
rect 1180 2395 1229 2407
rect 1180 1818 1188 2395
rect 1205 1818 1229 2395
rect 1180 1807 1229 1818
<< psubdiffcont >>
rect 414 1116 431 1191
rect 764 1116 781 1191
<< nsubdiffcont >>
rect -70 1822 -44 2392
rect 1188 1818 1205 2395
<< poly >>
rect 400 2485 751 2488
rect -90 2465 751 2485
rect 15 2406 65 2419
rect 115 2406 165 2419
rect 215 2406 265 2419
rect 401 2407 451 2465
rect 501 2407 551 2465
rect 601 2407 651 2465
rect 701 2407 751 2465
rect 880 2407 930 2422
rect 980 2407 1030 2422
rect 1080 2407 1130 2422
rect 15 1781 65 1806
rect 15 1756 23 1781
rect 55 1756 65 1781
rect 15 1751 65 1756
rect 115 1771 165 1806
rect 215 1771 265 1806
rect 401 1792 451 1807
rect 501 1792 551 1807
rect 601 1792 651 1807
rect 701 1792 751 1807
rect 880 1771 930 1807
rect 980 1771 1030 1807
rect 115 1736 1030 1771
rect 1080 1782 1130 1807
rect 1080 1747 1090 1782
rect 1120 1747 1130 1782
rect 1080 1742 1130 1747
rect 115 1730 140 1736
rect -90 1710 140 1730
rect -90 1666 235 1668
rect 401 1666 451 1667
rect -90 1646 550 1666
rect 181 1640 550 1646
rect -25 1616 130 1625
rect -25 1610 131 1616
rect -25 1606 10 1610
rect -25 1583 -17 1606
rect 2 1583 10 1606
rect 81 1602 131 1610
rect 181 1602 231 1640
rect 281 1602 351 1640
rect 401 1602 451 1640
rect 500 1616 550 1640
rect 500 1610 551 1616
rect 501 1602 551 1610
rect 601 1602 651 1615
rect 701 1602 751 1615
rect 801 1602 861 1615
rect 911 1602 961 1615
rect 1011 1602 1061 1615
rect -25 1575 10 1583
rect 81 1286 131 1301
rect 181 1286 231 1301
rect 281 1286 351 1301
rect 401 1286 451 1301
rect 501 1286 551 1301
rect 601 1286 651 1301
rect 701 1286 751 1301
rect 801 1286 861 1301
rect 601 1265 650 1286
rect 701 1265 750 1286
rect 801 1265 860 1286
rect 911 1265 961 1301
rect 1011 1286 1061 1301
rect 321 1264 961 1265
rect 21 1263 961 1264
rect -90 1240 961 1263
rect 1010 1260 1115 1286
rect -90 1239 960 1240
rect -90 1238 391 1239
rect -90 1237 196 1238
rect 115 1105 165 1115
rect -25 1090 16 1100
rect -25 1070 -15 1090
rect 4 1080 16 1090
rect 4 1070 65 1080
rect -25 1063 65 1070
rect 15 1050 65 1063
rect 115 1070 125 1105
rect 155 1070 165 1105
rect 115 1050 165 1070
rect 215 1050 265 1063
rect 401 1051 451 1064
rect 501 1051 551 1064
rect 601 1051 651 1064
rect 701 1051 751 1064
rect 880 1051 930 1066
rect 980 1051 1030 1066
rect 1080 1065 1115 1260
rect 1145 1220 1190 1230
rect 1145 1190 1155 1220
rect 1180 1195 1255 1220
rect 1180 1190 1190 1195
rect 1145 1180 1190 1190
rect 1080 1051 1130 1065
rect 15 435 65 450
rect 115 440 165 450
rect 215 440 265 450
rect 401 440 451 451
rect 501 440 551 451
rect 601 440 651 451
rect 701 440 751 451
rect 880 440 930 451
rect 980 440 1030 451
rect 115 431 1030 440
rect 115 425 990 431
rect 115 405 165 425
rect -90 382 165 405
rect 980 396 990 425
rect 1020 396 1030 431
rect 980 386 1030 396
rect -90 286 1030 308
rect 15 250 65 263
rect 115 250 165 286
rect 215 250 265 286
rect 401 251 451 264
rect 501 251 551 264
rect 601 251 651 264
rect 701 251 751 264
rect 880 251 930 286
rect 980 251 1030 286
rect 1080 251 1130 451
rect 15 -375 65 -350
rect 115 -365 165 -350
rect 215 -365 265 -350
rect 401 -357 451 -349
rect 501 -357 551 -349
rect 601 -357 651 -349
rect 701 -357 751 -349
rect 400 -365 751 -357
rect 880 -362 930 -349
rect 980 -362 1030 -349
rect 15 -410 25 -375
rect 55 -410 65 -375
rect 310 -373 751 -365
rect 310 -397 319 -373
rect 337 -384 751 -373
rect 337 -397 345 -384
rect 400 -385 751 -384
rect 1080 -369 1130 -349
rect 310 -403 345 -397
rect 1080 -404 1090 -369
rect 1120 -404 1130 -369
rect 1080 -409 1130 -404
rect 15 -417 65 -410
<< polycont >>
rect 23 1756 55 1781
rect 1090 1747 1120 1782
rect -17 1583 2 1606
rect -15 1070 4 1090
rect 125 1070 155 1105
rect 1155 1190 1180 1220
rect 990 396 1020 431
rect 25 -410 55 -375
rect 319 -397 337 -373
rect 1090 -404 1120 -369
<< locali >>
rect 70 2431 310 2451
rect -77 2396 10 2401
rect -77 2392 -20 2396
rect -77 1822 -70 2392
rect -44 1822 -20 2392
rect -77 1821 -20 1822
rect 0 1821 10 2396
rect -77 1811 10 1821
rect 70 2396 110 2431
rect 70 1821 80 2396
rect 100 1821 110 2396
rect 169 2396 210 2400
rect 169 2379 180 2396
rect 70 1811 110 1821
rect 170 1821 180 2379
rect 200 1821 210 2396
rect 15 1781 65 1792
rect 15 1756 23 1781
rect 55 1756 65 1781
rect 15 1751 65 1756
rect 170 1728 210 1821
rect 270 2396 310 2431
rect 835 2426 1076 2451
rect 270 1821 280 2396
rect 300 1821 310 2396
rect 270 1776 310 1821
rect 356 2397 396 2400
rect 356 1822 366 2397
rect 386 1822 396 2397
rect 356 1812 396 1822
rect 456 2397 496 2400
rect 456 1822 466 2397
rect 486 1822 496 2397
rect 456 1812 496 1822
rect 556 2397 596 2401
rect 556 1822 566 2397
rect 586 1822 596 2397
rect 556 1812 596 1822
rect 656 2397 696 2402
rect 656 1822 666 2397
rect 686 1822 696 2397
rect 656 1812 696 1822
rect 756 2397 796 2402
rect 756 1822 766 2397
rect 787 1822 796 2397
rect 756 1812 796 1822
rect 835 2392 875 2426
rect 835 1817 845 2392
rect 865 1817 875 2392
rect 356 1807 395 1812
rect 456 1776 495 1812
rect 556 1807 595 1812
rect 656 1790 695 1812
rect 756 1807 795 1812
rect 270 1749 495 1776
rect -55 1726 211 1728
rect -67 1687 211 1726
rect -67 376 -42 1687
rect 455 1652 495 1749
rect 235 1626 495 1652
rect -25 1606 10 1615
rect -25 1583 -17 1606
rect 2 1583 10 1606
rect 235 1602 275 1626
rect 456 1602 495 1626
rect 655 1776 695 1790
rect 835 1776 875 1817
rect 935 2392 975 2400
rect 935 1817 945 2392
rect 965 1834 975 2392
rect 1035 2393 1076 2426
rect 1135 2395 1214 2402
rect 1035 2392 1075 2393
rect 965 1817 976 1834
rect 935 1814 976 1817
rect 655 1751 875 1776
rect 655 1651 695 1751
rect 936 1716 976 1814
rect 1035 1817 1045 2392
rect 1065 1817 1075 2392
rect 1035 1807 1075 1817
rect 1135 2392 1188 2395
rect 1135 1817 1145 2392
rect 1165 1818 1188 2392
rect 1205 1818 1214 2395
rect 1165 1817 1214 1818
rect 1135 1812 1214 1817
rect 1080 1782 1130 1789
rect 1080 1747 1090 1782
rect 1120 1747 1130 1782
rect 1080 1742 1130 1747
rect 935 1691 1210 1716
rect 655 1625 905 1651
rect 565 1602 587 1603
rect 655 1602 695 1625
rect 865 1602 905 1625
rect -25 1575 10 1583
rect 36 1598 76 1602
rect 36 1316 46 1598
rect 66 1316 76 1598
rect 36 1313 76 1316
rect 136 1597 176 1602
rect 136 1316 146 1597
rect 166 1316 176 1597
rect 235 1598 276 1602
rect 235 1590 246 1598
rect 136 1306 176 1316
rect 236 1316 246 1590
rect 266 1316 276 1598
rect 236 1308 276 1316
rect 356 1597 396 1602
rect 356 1316 366 1597
rect 386 1316 396 1597
rect 356 1306 396 1316
rect 136 1265 175 1306
rect 355 1265 396 1306
rect 456 1598 496 1602
rect 456 1316 466 1598
rect 486 1316 496 1598
rect 556 1598 596 1602
rect 556 1316 566 1598
rect 586 1316 596 1598
rect 655 1597 696 1602
rect 655 1590 666 1597
rect 456 1306 496 1316
rect 456 1301 495 1306
rect 555 1265 596 1316
rect 656 1316 666 1590
rect 686 1316 696 1597
rect 656 1306 696 1316
rect 756 1597 794 1602
rect 756 1316 766 1597
rect 786 1316 794 1597
rect 865 1597 906 1602
rect 865 1592 876 1597
rect 656 1301 695 1306
rect 756 1265 794 1316
rect 866 1316 876 1592
rect 896 1316 906 1597
rect 866 1308 906 1316
rect 966 1597 1006 1602
rect 966 1316 976 1597
rect 996 1316 1006 1597
rect 966 1314 1006 1316
rect 965 1308 1006 1314
rect 1066 1597 1106 1602
rect 1066 1315 1076 1597
rect 1096 1315 1106 1597
rect 1066 1309 1106 1315
rect 965 1265 1005 1308
rect 136 1250 1005 1265
rect 136 1240 1001 1250
rect 404 1191 442 1200
rect 404 1116 414 1191
rect 431 1116 442 1191
rect 115 1105 165 1115
rect 404 1106 442 1116
rect 115 1101 125 1105
rect -25 1090 16 1100
rect -25 1070 -15 1090
rect 4 1070 16 1090
rect -25 1063 16 1070
rect 78 1075 125 1101
rect 78 1045 96 1075
rect 115 1070 125 1075
rect 155 1070 165 1105
rect 115 1063 165 1070
rect -25 1035 10 1045
rect -25 470 -15 1035
rect 2 470 10 1035
rect -25 455 10 470
rect 70 1040 110 1045
rect 70 465 80 1040
rect 100 465 110 1040
rect 169 1040 210 1044
rect 169 1023 180 1040
rect 70 425 110 465
rect 170 465 180 1023
rect 200 465 210 1040
rect 170 455 210 465
rect 270 1040 310 1045
rect 270 465 280 1040
rect 300 465 310 1040
rect 270 425 310 465
rect 356 1041 396 1051
rect 356 466 366 1041
rect 386 466 396 1041
rect 356 458 396 466
rect 70 398 310 425
rect 355 456 396 458
rect 456 1046 495 1049
rect 456 1041 496 1046
rect 456 466 465 1041
rect 486 466 496 1041
rect 555 1045 594 1240
rect 1190 1230 1210 1691
rect 1145 1220 1210 1230
rect 754 1191 792 1200
rect 754 1116 764 1191
rect 781 1116 792 1191
rect 1145 1190 1155 1220
rect 1180 1190 1210 1220
rect 1145 1180 1210 1190
rect 754 1106 792 1116
rect 835 1076 1075 1103
rect 555 1041 596 1045
rect 555 1040 566 1041
rect 556 466 566 1040
rect 586 466 596 1041
rect 456 456 496 466
rect 355 430 395 456
rect 456 451 495 456
rect 555 430 596 466
rect 656 1041 696 1046
rect 656 466 666 1041
rect 686 466 696 1041
rect 656 458 696 466
rect 756 1041 796 1046
rect 756 466 766 1041
rect 786 466 796 1041
rect 756 456 796 466
rect 835 1036 875 1076
rect 835 461 845 1036
rect 865 461 875 1036
rect 835 456 875 461
rect 935 1036 975 1046
rect 1034 1042 1075 1076
rect 935 461 945 1036
rect 965 478 975 1036
rect 1035 1036 1075 1042
rect 965 461 976 478
rect 935 457 976 461
rect 1035 461 1045 1036
rect 1065 461 1075 1036
rect 1035 456 1075 461
rect 1135 1036 1172 1046
rect 1135 461 1143 1036
rect 1163 461 1172 1036
rect 1135 456 1172 461
rect 756 430 795 456
rect 355 410 795 430
rect 980 431 1030 438
rect 980 396 990 431
rect 1020 430 1030 431
rect 1050 430 1075 456
rect 1020 400 1075 430
rect 1020 396 1030 400
rect 980 386 1030 396
rect -67 355 105 376
rect 1190 365 1210 1180
rect 82 245 105 355
rect 170 282 495 307
rect 1189 305 1210 365
rect 170 250 210 282
rect -30 240 10 245
rect -30 -335 -20 240
rect 1 -335 10 240
rect -30 -345 10 -335
rect 70 240 110 245
rect 70 -335 80 240
rect 100 -335 110 240
rect 169 240 210 250
rect 169 223 180 240
rect 70 -338 110 -335
rect 82 -341 110 -338
rect 170 -335 180 223
rect 200 -335 210 240
rect 15 -375 65 -365
rect 15 -410 25 -375
rect 55 -410 65 -375
rect 82 -375 111 -341
rect 170 -345 210 -335
rect 270 240 310 245
rect 270 -335 280 240
rect 300 -335 310 240
rect 270 -365 310 -335
rect 356 242 396 251
rect 356 -333 365 242
rect 356 -334 366 -333
rect 386 -334 396 242
rect 455 246 495 282
rect 835 278 1210 305
rect 455 241 496 246
rect 455 240 466 241
rect 356 -344 396 -334
rect 456 -334 466 240
rect 486 -334 496 241
rect 456 -344 496 -334
rect 556 241 596 245
rect 556 -335 566 241
rect 586 240 596 241
rect 587 -335 596 240
rect 556 -344 596 -335
rect 656 241 696 246
rect 656 -334 666 241
rect 686 -334 696 241
rect 656 -344 696 -334
rect 756 241 796 246
rect 756 -335 766 241
rect 786 240 796 241
rect 787 -335 796 240
rect 756 -344 796 -335
rect 835 236 875 278
rect 835 -339 845 236
rect 865 -339 875 236
rect 835 -344 875 -339
rect 935 236 975 246
rect 1034 242 1075 278
rect 935 -339 945 236
rect 965 -322 975 236
rect 1035 236 1075 242
rect 965 -339 976 -322
rect 356 -349 395 -344
rect 456 -349 495 -344
rect 556 -349 595 -344
rect 270 -373 345 -365
rect 270 -375 319 -373
rect 82 -397 319 -375
rect 337 -397 345 -373
rect 82 -402 345 -397
rect 656 -375 695 -344
rect 756 -349 795 -344
rect 935 -349 976 -339
rect 1035 -339 1045 236
rect 1065 -339 1075 236
rect 1035 -344 1075 -339
rect 1135 236 1175 246
rect 1135 -339 1145 236
rect 1166 -339 1175 236
rect 1135 -344 1175 -339
rect 935 -375 975 -349
rect 656 -400 975 -375
rect 1080 -369 1130 -362
rect 310 -403 345 -402
rect 1080 -404 1090 -369
rect 1120 -404 1130 -369
rect 1080 -409 1130 -404
rect 15 -417 65 -410
<< viali >>
rect -70 1822 -44 2392
rect -20 1821 0 2396
rect 23 1756 55 1781
rect 366 1822 386 2397
rect 566 1822 586 2397
rect 767 1822 786 2397
rect 786 1822 787 2397
rect -17 1583 2 1606
rect 1145 1817 1165 2392
rect 1188 1818 1205 2395
rect 1090 1747 1120 1782
rect 46 1316 66 1598
rect 1076 1316 1096 1597
rect 1076 1315 1096 1316
rect 414 1116 431 1191
rect -15 1070 4 1090
rect -15 470 2 1035
rect 180 465 200 1040
rect 465 466 466 1041
rect 466 466 485 1041
rect 764 1116 781 1191
rect 666 466 686 1041
rect 945 461 965 1036
rect 1143 461 1163 1036
rect -20 -335 0 240
rect 0 -335 1 240
rect 25 -410 55 -375
rect 365 241 386 242
rect 365 -333 366 241
rect 366 -333 386 241
rect 566 -334 586 240
rect 586 -334 587 240
rect 566 -335 587 -334
rect 766 -334 786 240
rect 786 -334 787 240
rect 766 -335 787 -334
rect 1145 -339 1165 236
rect 1165 -339 1166 236
rect 1090 -404 1120 -369
<< metal1 >>
rect -58 2443 1208 2458
rect -94 2397 1250 2443
rect -94 2396 366 2397
rect -94 2392 -20 2396
rect -94 1822 -70 2392
rect -44 1822 -20 2392
rect -94 1821 -20 1822
rect 0 1822 366 2396
rect 386 1822 566 2397
rect 586 1822 767 2397
rect 787 2395 1250 2397
rect 787 2392 1188 2395
rect 787 1822 1145 2392
rect 0 1821 1145 1822
rect -94 1817 1145 1821
rect 1165 1818 1188 2392
rect 1205 1818 1250 2395
rect 1165 1817 1250 1818
rect -94 1792 1250 1817
rect -94 1791 1208 1792
rect -58 1782 1208 1791
rect -58 1781 1090 1782
rect -58 1756 23 1781
rect 55 1756 1090 1781
rect -58 1747 1090 1756
rect 1120 1747 1208 1782
rect -58 1722 1208 1747
rect -60 1606 1196 1671
rect -60 1583 -17 1606
rect 2 1598 1196 1606
rect 2 1583 46 1598
rect -60 1316 46 1583
rect 66 1597 1196 1598
rect 66 1316 1076 1597
rect -60 1315 1076 1316
rect 1096 1315 1196 1597
rect -60 1191 1196 1315
rect -60 1116 414 1191
rect 431 1116 764 1191
rect 781 1116 1196 1191
rect -60 1090 1196 1116
rect -60 1070 -15 1090
rect 4 1070 1196 1090
rect -60 1041 1196 1070
rect -60 1040 465 1041
rect -60 1035 180 1040
rect -60 470 -15 1035
rect 2 470 180 1035
rect -60 465 180 470
rect 200 466 465 1040
rect 485 466 666 1041
rect 686 1036 1196 1041
rect 686 466 945 1036
rect 200 465 945 466
rect -60 461 945 465
rect 965 461 1143 1036
rect 1163 461 1196 1036
rect -60 242 1196 461
rect -60 240 365 242
rect -60 -335 -20 240
rect 1 -333 365 240
rect 386 240 1196 242
rect 386 -333 566 240
rect 1 -335 566 -333
rect 587 -335 766 240
rect 787 236 1196 240
rect 787 -335 1145 236
rect -60 -339 1145 -335
rect 1166 -339 1196 236
rect -60 -369 1196 -339
rect -60 -375 1090 -369
rect -60 -410 25 -375
rect 55 -404 1090 -375
rect 1120 -404 1196 -369
rect 55 -410 1196 -404
rect -60 -434 1196 -410
<< labels >>
rlabel poly -90 1655 -90 1655 7 V1
rlabel poly -90 1720 -90 1720 7 Vcp
rlabel metal1 -58 2455 -58 2455 7 Vp
rlabel poly -90 2475 -90 2475 7 Vbp
rlabel poly -90 1250 -90 1250 7 V2
rlabel poly 1255 1205 1255 1205 3 Vout
rlabel poly -90 392 -90 392 3 Vbn
rlabel poly -90 294 -90 294 3 Vcn
rlabel metal1 -60 330 -60 330 7 VN
<< end >>
