magic
tech sky130A
timestamp 1697386427
<< nwell >>
rect -68 2495 1201 2496
rect -90 1716 1257 2495
<< nmos >>
rect 81 1001 131 1601
rect 181 1001 231 1601
rect 281 1001 351 1601
rect 401 1001 451 1601
rect 501 1001 551 1601
rect 601 1001 651 1601
rect 701 1001 751 1601
rect 801 1001 861 1601
rect 911 1001 961 1601
rect 1011 1001 1061 1601
rect 15 200 65 800
rect 115 200 165 800
rect 215 200 265 800
rect 401 201 451 801
rect 501 201 551 801
rect 601 201 651 801
rect 701 201 751 801
rect 880 201 930 801
rect 980 201 1030 801
rect 1080 201 1130 801
rect 15 -600 65 0
rect 115 -600 165 0
rect 215 -600 265 0
rect 401 -599 451 1
rect 501 -599 551 1
rect 601 -599 651 1
rect 701 -599 751 1
rect 880 -599 930 1
rect 980 -599 1030 1
rect 1080 -599 1130 1
<< pmos >>
rect 15 1806 65 2406
rect 115 1806 165 2406
rect 215 1806 265 2406
rect 401 1807 451 2407
rect 501 1807 551 2407
rect 601 1807 651 2407
rect 701 1807 751 2407
rect 880 1807 930 2407
rect 980 1807 1030 2407
rect 1080 1807 1130 2407
<< ndiff >>
rect 31 1591 81 1601
rect 31 1016 46 1591
rect 66 1016 81 1591
rect 31 1001 81 1016
rect 131 1591 181 1601
rect 131 1016 146 1591
rect 166 1016 181 1591
rect 131 1001 181 1016
rect 231 1591 281 1601
rect 231 1016 246 1591
rect 266 1016 281 1591
rect 231 1001 281 1016
rect 351 1591 401 1601
rect 351 1016 366 1591
rect 386 1016 401 1591
rect 351 1001 401 1016
rect 451 1591 501 1601
rect 451 1016 466 1591
rect 486 1016 501 1591
rect 451 1001 501 1016
rect 551 1591 601 1601
rect 551 1016 566 1591
rect 586 1016 601 1591
rect 551 1001 601 1016
rect 651 1591 701 1601
rect 651 1016 666 1591
rect 686 1016 701 1591
rect 651 1001 701 1016
rect 751 1591 801 1601
rect 751 1016 766 1591
rect 786 1016 801 1591
rect 751 1001 801 1016
rect 861 1591 911 1601
rect 861 1016 876 1591
rect 896 1016 911 1591
rect 861 1001 911 1016
rect 961 1591 1011 1601
rect 961 1016 976 1591
rect 996 1016 1011 1591
rect 961 1001 1011 1016
rect 1061 1591 1109 1601
rect 1061 1016 1076 1591
rect 1096 1016 1109 1591
rect 1061 1001 1109 1016
rect -35 785 15 800
rect -35 220 -15 785
rect 2 220 15 785
rect -35 200 15 220
rect 65 790 115 800
rect 65 215 80 790
rect 100 215 115 790
rect 65 200 115 215
rect 165 790 215 800
rect 165 215 180 790
rect 200 215 215 790
rect 165 200 215 215
rect 265 790 315 800
rect 265 215 280 790
rect 300 215 315 790
rect 265 200 315 215
rect 351 791 401 801
rect 351 216 366 791
rect 386 216 401 791
rect 351 201 401 216
rect 451 791 501 801
rect 451 216 466 791
rect 486 216 501 791
rect 451 201 501 216
rect 551 791 601 801
rect 551 216 566 791
rect 586 216 601 791
rect 551 201 601 216
rect 651 791 701 801
rect 651 216 666 791
rect 686 216 701 791
rect 651 201 701 216
rect 751 791 799 801
rect 751 216 766 791
rect 786 216 799 791
rect 751 201 799 216
rect 830 786 880 801
rect 830 211 845 786
rect 865 211 880 786
rect 830 201 880 211
rect 930 786 980 801
rect 930 211 945 786
rect 965 211 980 786
rect 930 201 980 211
rect 1030 786 1080 801
rect 1030 211 1045 786
rect 1065 211 1080 786
rect 1030 201 1080 211
rect 1130 786 1180 801
rect 1130 211 1143 786
rect 1163 211 1180 786
rect 1130 201 1180 211
rect -35 -10 15 0
rect -35 -585 -20 -10
rect 0 -585 15 -10
rect -35 -600 15 -585
rect 65 -10 115 0
rect 65 -585 80 -10
rect 100 -585 115 -10
rect 65 -600 115 -585
rect 165 -10 215 0
rect 165 -585 180 -10
rect 200 -585 215 -10
rect 165 -600 215 -585
rect 265 -10 315 0
rect 265 -585 280 -10
rect 300 -585 315 -10
rect 265 -600 315 -585
rect 351 -9 401 1
rect 351 -584 366 -9
rect 386 -584 401 -9
rect 351 -599 401 -584
rect 451 -9 501 1
rect 451 -584 466 -9
rect 486 -584 501 -9
rect 451 -599 501 -584
rect 551 -9 601 1
rect 551 -584 566 -9
rect 586 -584 601 -9
rect 551 -599 601 -584
rect 651 -9 701 1
rect 651 -584 666 -9
rect 686 -584 701 -9
rect 651 -599 701 -584
rect 751 -9 799 1
rect 751 -584 766 -9
rect 786 -584 799 -9
rect 751 -599 799 -584
rect 830 -14 880 1
rect 830 -589 845 -14
rect 865 -589 880 -14
rect 830 -599 880 -589
rect 930 -14 980 1
rect 930 -589 945 -14
rect 965 -589 980 -14
rect 930 -599 980 -589
rect 1030 -14 1080 1
rect 1030 -589 1045 -14
rect 1065 -589 1080 -14
rect 1030 -599 1080 -589
rect 1130 -14 1180 1
rect 1130 -589 1145 -14
rect 1165 -589 1180 -14
rect 1130 -599 1180 -589
<< pdiff >>
rect -35 2396 15 2406
rect -35 1821 -20 2396
rect 0 1821 15 2396
rect -35 1806 15 1821
rect 65 2396 115 2406
rect 65 1821 80 2396
rect 100 1821 115 2396
rect 65 1806 115 1821
rect 165 2396 215 2406
rect 165 1821 180 2396
rect 200 1821 215 2396
rect 165 1806 215 1821
rect 265 2396 315 2406
rect 265 1821 280 2396
rect 300 1821 315 2396
rect 265 1806 315 1821
rect 351 2397 401 2407
rect 351 1822 366 2397
rect 386 1822 401 2397
rect 351 1807 401 1822
rect 451 2397 501 2407
rect 451 1822 466 2397
rect 486 1822 501 2397
rect 451 1807 501 1822
rect 551 2397 601 2407
rect 551 1822 566 2397
rect 586 1822 601 2397
rect 551 1807 601 1822
rect 651 2397 701 2407
rect 651 1822 666 2397
rect 686 1822 701 2397
rect 651 1807 701 1822
rect 751 2397 799 2407
rect 751 1822 766 2397
rect 786 1822 799 2397
rect 751 1807 799 1822
rect 830 2392 880 2407
rect 830 1817 845 2392
rect 865 1817 880 2392
rect 830 1807 880 1817
rect 930 2392 980 2407
rect 930 1817 945 2392
rect 965 1817 980 2392
rect 930 1807 980 1817
rect 1030 2392 1080 2407
rect 1030 1817 1045 2392
rect 1065 1817 1080 2392
rect 1030 1807 1080 1817
rect 1130 2392 1180 2407
rect 1130 1817 1145 2392
rect 1165 1817 1180 2392
rect 1130 1807 1180 1817
<< ndiffc >>
rect 46 1016 66 1591
rect 146 1016 166 1591
rect 246 1016 266 1591
rect 366 1016 386 1591
rect 466 1016 486 1591
rect 566 1016 586 1591
rect 666 1016 686 1591
rect 766 1016 786 1591
rect 876 1016 896 1591
rect 976 1016 996 1591
rect 1076 1016 1096 1591
rect -15 220 2 785
rect 80 215 100 790
rect 180 215 200 790
rect 280 215 300 790
rect 366 216 386 791
rect 466 216 486 791
rect 566 216 586 791
rect 666 216 686 791
rect 766 216 786 791
rect 845 211 865 786
rect 945 211 965 786
rect 1045 211 1065 786
rect 1143 211 1163 786
rect -20 -585 0 -10
rect 80 -585 100 -10
rect 180 -585 200 -10
rect 280 -585 300 -10
rect 366 -584 386 -9
rect 466 -584 486 -9
rect 566 -584 586 -9
rect 666 -584 686 -9
rect 766 -584 786 -9
rect 845 -589 865 -14
rect 945 -589 965 -14
rect 1045 -589 1065 -14
rect 1145 -589 1165 -14
<< pdiffc >>
rect -20 1821 0 2396
rect 80 1821 100 2396
rect 180 1821 200 2396
rect 280 1821 300 2396
rect 366 1822 386 2397
rect 466 1822 486 2397
rect 566 1822 586 2397
rect 666 1822 686 2397
rect 766 1822 786 2397
rect 845 1817 865 2392
rect 945 1817 965 2392
rect 1045 1817 1065 2392
rect 1145 1817 1165 2392
<< poly >>
rect 400 2485 751 2488
rect -90 2465 751 2485
rect 15 2406 65 2419
rect 115 2406 165 2419
rect 215 2406 265 2419
rect 401 2407 451 2465
rect 501 2407 551 2465
rect 601 2407 651 2465
rect 701 2407 751 2465
rect 880 2407 930 2422
rect 980 2407 1030 2422
rect 1080 2407 1130 2422
rect 15 1781 65 1806
rect 15 1756 23 1781
rect 55 1756 65 1781
rect 15 1751 65 1756
rect 115 1771 165 1806
rect 215 1771 265 1806
rect 401 1792 451 1807
rect 501 1792 551 1807
rect 601 1792 651 1807
rect 701 1792 751 1807
rect 880 1771 930 1807
rect 980 1771 1030 1807
rect 115 1736 1030 1771
rect 1080 1782 1130 1807
rect 1080 1747 1090 1782
rect 1120 1747 1130 1782
rect 1080 1742 1130 1747
rect 115 1730 140 1736
rect -90 1710 140 1730
rect -90 1666 235 1668
rect 401 1666 451 1667
rect -90 1646 550 1666
rect 181 1640 550 1646
rect -25 1616 130 1625
rect -25 1609 131 1616
rect -25 1606 10 1609
rect -25 1583 -17 1606
rect 2 1583 10 1606
rect 81 1601 131 1609
rect 181 1601 231 1640
rect 281 1601 351 1640
rect 401 1601 451 1640
rect 500 1614 550 1640
rect 500 1610 551 1614
rect 501 1601 551 1610
rect 601 1601 651 1614
rect 701 1601 751 1614
rect 801 1601 861 1614
rect 911 1601 961 1614
rect 1011 1601 1061 1614
rect -25 1575 10 1583
rect 81 986 131 1001
rect 181 986 231 1001
rect 281 986 351 1001
rect 401 986 451 1001
rect 501 986 551 1001
rect 601 986 651 1001
rect 701 986 751 1001
rect 801 986 861 1001
rect 601 965 650 986
rect 701 965 750 986
rect 801 965 860 986
rect 911 965 961 1001
rect 1011 986 1061 1001
rect 321 964 961 965
rect 21 963 961 964
rect -90 940 961 963
rect 1010 960 1115 986
rect -90 939 960 940
rect -90 938 391 939
rect -90 937 196 938
rect 115 855 165 865
rect -25 840 16 850
rect -25 820 -15 840
rect 4 830 16 840
rect 4 820 65 830
rect -25 813 65 820
rect 15 800 65 813
rect 115 820 125 855
rect 155 820 165 855
rect 115 800 165 820
rect 215 800 265 813
rect 401 801 451 814
rect 501 801 551 814
rect 601 801 651 814
rect 701 801 751 814
rect 880 801 930 816
rect 980 801 1030 816
rect 1080 815 1115 960
rect 1145 920 1190 930
rect 1145 890 1155 920
rect 1180 895 1255 920
rect 1180 890 1190 895
rect 1145 880 1190 890
rect 1080 801 1130 815
rect 15 185 65 200
rect 115 190 165 200
rect 215 190 265 200
rect 401 190 451 201
rect 501 190 551 201
rect 601 190 651 201
rect 701 190 751 201
rect 880 190 930 201
rect 980 190 1030 201
rect 115 181 1030 190
rect 115 175 990 181
rect 115 155 165 175
rect -90 132 165 155
rect 980 146 990 175
rect 1020 146 1030 181
rect 980 136 1030 146
rect -90 36 1030 58
rect 15 0 65 13
rect 115 0 165 36
rect 215 0 265 36
rect 401 1 451 14
rect 501 1 551 14
rect 601 1 651 14
rect 701 1 751 14
rect 880 1 930 36
rect 980 1 1030 36
rect 1080 1 1130 201
rect 15 -625 65 -600
rect 115 -615 165 -600
rect 215 -615 265 -600
rect 401 -607 451 -599
rect 501 -607 551 -599
rect 601 -607 651 -599
rect 701 -607 751 -599
rect 400 -615 751 -607
rect 880 -612 930 -599
rect 980 -612 1030 -599
rect 15 -660 25 -625
rect 55 -660 65 -625
rect 310 -623 751 -615
rect 310 -647 319 -623
rect 337 -634 751 -623
rect 337 -647 345 -634
rect 400 -635 751 -634
rect 1080 -619 1130 -599
rect 310 -653 345 -647
rect 1080 -654 1090 -619
rect 1120 -654 1130 -619
rect 1080 -659 1130 -654
rect 15 -667 65 -660
<< polycont >>
rect 23 1756 55 1781
rect 1090 1747 1120 1782
rect -17 1583 2 1606
rect -15 820 4 840
rect 125 820 155 855
rect 1155 890 1180 920
rect 990 146 1020 181
rect 25 -660 55 -625
rect 319 -647 337 -623
rect 1090 -654 1120 -619
<< locali >>
rect 70 2431 310 2451
rect -30 2396 10 2401
rect -30 1821 -20 2396
rect 0 1821 10 2396
rect -30 1811 10 1821
rect 70 2396 110 2431
rect 70 1821 80 2396
rect 100 1821 110 2396
rect 169 2396 210 2400
rect 169 2379 180 2396
rect 70 1811 110 1821
rect 170 1821 180 2379
rect 200 1821 210 2396
rect 15 1781 65 1792
rect 15 1756 23 1781
rect 55 1756 65 1781
rect 15 1751 65 1756
rect 170 1728 210 1821
rect 270 2396 310 2431
rect 835 2426 1076 2451
rect 270 1821 280 2396
rect 300 1821 310 2396
rect 270 1776 310 1821
rect 356 2397 396 2400
rect 356 1822 366 2397
rect 386 1822 396 2397
rect 356 1812 396 1822
rect 456 2397 496 2400
rect 456 1822 466 2397
rect 486 1822 496 2397
rect 456 1812 496 1822
rect 556 2397 596 2401
rect 556 1822 566 2397
rect 586 1822 596 2397
rect 556 1812 596 1822
rect 656 2397 696 2402
rect 656 1822 666 2397
rect 686 1822 696 2397
rect 656 1812 696 1822
rect 756 2397 796 2402
rect 756 1822 766 2397
rect 787 1822 796 2397
rect 756 1812 796 1822
rect 835 2392 875 2426
rect 835 1817 845 2392
rect 865 1817 875 2392
rect 356 1807 395 1812
rect 456 1776 495 1812
rect 556 1807 595 1812
rect 656 1790 695 1812
rect 756 1807 795 1812
rect 270 1749 495 1776
rect -55 1726 211 1728
rect -67 1687 211 1726
rect -67 126 -42 1687
rect 455 1652 495 1749
rect 235 1626 495 1652
rect -25 1606 10 1615
rect -25 1583 -17 1606
rect 2 1583 10 1606
rect 235 1601 275 1626
rect -25 1575 10 1583
rect 36 1592 76 1595
rect 36 1016 46 1592
rect 66 1016 76 1592
rect 36 1013 76 1016
rect 136 1591 176 1595
rect 136 1016 146 1591
rect 166 1016 176 1591
rect 235 1591 276 1601
rect 456 1596 495 1626
rect 655 1776 695 1790
rect 835 1776 875 1817
rect 935 2392 975 2400
rect 935 1817 945 2392
rect 965 1834 975 2392
rect 1035 2393 1076 2426
rect 1035 2392 1075 2393
rect 965 1817 976 1834
rect 935 1814 976 1817
rect 655 1751 875 1776
rect 655 1651 695 1751
rect 936 1716 976 1814
rect 1035 1817 1045 2392
rect 1065 1817 1075 2392
rect 1035 1807 1075 1817
rect 1135 2392 1175 2402
rect 1135 1817 1145 2392
rect 1165 1817 1175 2392
rect 1135 1812 1175 1817
rect 1080 1782 1130 1789
rect 1080 1747 1090 1782
rect 1120 1747 1130 1782
rect 1080 1742 1130 1747
rect 935 1691 1210 1716
rect 655 1625 905 1651
rect 655 1601 695 1625
rect 235 1590 246 1591
rect 136 1006 176 1016
rect 236 1016 246 1590
rect 266 1016 276 1591
rect 236 1008 276 1016
rect 356 1591 396 1595
rect 356 1016 366 1591
rect 386 1016 396 1591
rect 356 1006 396 1016
rect 136 965 175 1006
rect 355 965 396 1006
rect 456 1591 496 1596
rect 456 1016 466 1591
rect 486 1016 496 1591
rect 556 1591 596 1601
rect 556 1016 566 1591
rect 586 1016 596 1591
rect 655 1591 696 1601
rect 655 1590 666 1591
rect 456 1006 496 1016
rect 456 1001 495 1006
rect 555 965 596 1016
rect 656 1016 666 1590
rect 686 1016 696 1591
rect 656 1006 696 1016
rect 756 1591 794 1599
rect 865 1596 905 1625
rect 865 1592 906 1596
rect 756 1016 766 1591
rect 786 1016 794 1591
rect 656 1001 695 1006
rect 756 965 794 1016
rect 866 1591 906 1592
rect 866 1016 876 1591
rect 896 1016 906 1591
rect 866 1008 906 1016
rect 966 1591 1006 1596
rect 966 1016 976 1591
rect 996 1016 1006 1591
rect 966 1014 1006 1016
rect 965 1008 1006 1014
rect 1066 1591 1106 1596
rect 1066 1015 1076 1591
rect 1096 1015 1106 1591
rect 1066 1009 1106 1015
rect 965 965 1005 1008
rect 136 950 1005 965
rect 136 940 1001 950
rect 115 855 165 865
rect 115 851 125 855
rect -25 840 16 850
rect -25 820 -15 840
rect 4 820 16 840
rect -25 813 16 820
rect 78 825 125 851
rect 78 795 96 825
rect 115 820 125 825
rect 155 820 165 855
rect 115 813 165 820
rect -25 785 10 795
rect -25 220 -15 785
rect 2 220 10 785
rect -25 205 10 220
rect 70 790 110 795
rect 70 215 80 790
rect 100 215 110 790
rect 169 790 210 794
rect 169 773 180 790
rect 70 175 110 215
rect 170 215 180 773
rect 200 215 210 790
rect 170 205 210 215
rect 270 790 310 795
rect 270 215 280 790
rect 300 215 310 790
rect 270 175 310 215
rect 356 791 396 801
rect 356 216 366 791
rect 386 216 396 791
rect 356 208 396 216
rect 70 148 310 175
rect 355 206 396 208
rect 456 796 495 799
rect 456 791 496 796
rect 456 216 465 791
rect 486 216 496 791
rect 555 795 594 940
rect 1190 930 1210 1691
rect 1145 920 1210 930
rect 1145 890 1155 920
rect 1180 890 1210 920
rect 1145 880 1210 890
rect 835 826 1075 853
rect 555 791 596 795
rect 555 790 566 791
rect 556 216 566 790
rect 586 216 596 791
rect 456 206 496 216
rect 355 180 395 206
rect 456 201 495 206
rect 555 180 596 216
rect 656 791 696 796
rect 656 216 666 791
rect 686 216 696 791
rect 656 208 696 216
rect 756 791 796 796
rect 756 216 766 791
rect 786 216 796 791
rect 756 206 796 216
rect 835 786 875 826
rect 835 211 845 786
rect 865 211 875 786
rect 835 206 875 211
rect 935 786 975 796
rect 1034 792 1075 826
rect 935 211 945 786
rect 965 228 975 786
rect 1035 786 1075 792
rect 965 211 976 228
rect 935 207 976 211
rect 1035 211 1045 786
rect 1065 211 1075 786
rect 1035 206 1075 211
rect 1135 786 1172 796
rect 1135 211 1143 786
rect 1163 211 1172 786
rect 1135 206 1172 211
rect 756 180 795 206
rect 355 160 795 180
rect 980 181 1030 188
rect 980 146 990 181
rect 1020 180 1030 181
rect 1050 180 1075 206
rect 1020 150 1075 180
rect 1020 146 1030 150
rect 980 136 1030 146
rect -67 105 105 126
rect 1190 115 1210 880
rect 82 -5 105 105
rect 170 32 495 57
rect 1189 55 1210 115
rect 170 0 210 32
rect -30 -10 10 -5
rect -30 -585 -20 -10
rect 1 -585 10 -10
rect -30 -595 10 -585
rect 70 -10 110 -5
rect 70 -585 80 -10
rect 100 -585 110 -10
rect 169 -10 210 0
rect 169 -27 180 -10
rect 70 -588 110 -585
rect 82 -591 110 -588
rect 170 -585 180 -27
rect 200 -585 210 -10
rect 15 -625 65 -615
rect 15 -660 25 -625
rect 55 -660 65 -625
rect 82 -625 111 -591
rect 170 -595 210 -585
rect 270 -10 310 -5
rect 270 -585 280 -10
rect 300 -585 310 -10
rect 270 -615 310 -585
rect 356 -8 396 1
rect 356 -583 365 -8
rect 356 -584 366 -583
rect 386 -584 396 -8
rect 455 -4 495 32
rect 835 28 1210 55
rect 455 -9 496 -4
rect 455 -10 466 -9
rect 356 -594 396 -584
rect 456 -584 466 -10
rect 486 -584 496 -9
rect 456 -594 496 -584
rect 556 -9 596 -5
rect 556 -585 566 -9
rect 586 -10 596 -9
rect 587 -585 596 -10
rect 556 -594 596 -585
rect 656 -9 696 -4
rect 656 -584 666 -9
rect 686 -584 696 -9
rect 656 -594 696 -584
rect 756 -9 796 -4
rect 756 -585 766 -9
rect 786 -10 796 -9
rect 787 -585 796 -10
rect 756 -594 796 -585
rect 835 -14 875 28
rect 835 -589 845 -14
rect 865 -589 875 -14
rect 835 -594 875 -589
rect 935 -14 975 -4
rect 1034 -8 1075 28
rect 935 -589 945 -14
rect 965 -572 975 -14
rect 1035 -14 1075 -8
rect 965 -589 976 -572
rect 356 -599 395 -594
rect 456 -599 495 -594
rect 556 -599 595 -594
rect 270 -623 345 -615
rect 270 -625 319 -623
rect 82 -647 319 -625
rect 337 -647 345 -623
rect 82 -652 345 -647
rect 656 -625 695 -594
rect 756 -599 795 -594
rect 935 -599 976 -589
rect 1035 -589 1045 -14
rect 1065 -589 1075 -14
rect 1035 -594 1075 -589
rect 1135 -14 1175 -4
rect 1135 -589 1145 -14
rect 1166 -589 1175 -14
rect 1135 -594 1175 -589
rect 935 -625 975 -599
rect 656 -650 975 -625
rect 1080 -619 1130 -612
rect 310 -653 345 -652
rect 1080 -654 1090 -619
rect 1120 -654 1130 -619
rect 1080 -659 1130 -654
rect 15 -667 65 -660
<< viali >>
rect -20 1821 0 2396
rect 23 1756 55 1781
rect 366 1822 386 2397
rect 566 1822 586 2397
rect 767 1822 786 2397
rect 786 1822 787 2397
rect -17 1583 2 1606
rect 46 1591 66 1592
rect 46 1016 66 1591
rect 1145 1817 1165 2392
rect 1090 1747 1120 1782
rect 1076 1016 1096 1591
rect 1076 1015 1096 1016
rect -15 820 4 840
rect -15 220 2 785
rect 180 215 200 790
rect 465 216 466 791
rect 466 216 485 791
rect 666 216 686 791
rect 945 211 965 786
rect 1143 211 1163 786
rect -20 -585 0 -10
rect 0 -585 1 -10
rect 25 -660 55 -625
rect 365 -9 386 -8
rect 365 -583 366 -9
rect 366 -583 386 -9
rect 566 -584 586 -10
rect 586 -584 587 -10
rect 566 -585 587 -584
rect 766 -584 786 -10
rect 786 -584 787 -10
rect 766 -585 787 -584
rect 1145 -589 1165 -14
rect 1165 -589 1166 -14
rect 1090 -654 1120 -619
<< metal1 >>
rect -58 2397 1208 2458
rect -58 2396 366 2397
rect -58 1821 -20 2396
rect 0 1822 366 2396
rect 386 1822 566 2397
rect 586 1822 767 2397
rect 787 2392 1208 2397
rect 787 1822 1145 2392
rect 0 1821 1145 1822
rect -58 1817 1145 1821
rect 1165 1817 1208 2392
rect -58 1782 1208 1817
rect -58 1781 1090 1782
rect -58 1756 23 1781
rect 55 1756 1090 1781
rect -58 1747 1090 1756
rect 1120 1747 1208 1782
rect -58 1722 1208 1747
rect -60 1606 1196 1671
rect -60 1583 -17 1606
rect 2 1592 1196 1606
rect 2 1583 46 1592
rect -60 1016 46 1583
rect 66 1591 1196 1592
rect 66 1016 1076 1591
rect -60 1015 1076 1016
rect 1096 1015 1196 1591
rect -60 840 1196 1015
rect -60 820 -15 840
rect 4 820 1196 840
rect -60 791 1196 820
rect -60 790 465 791
rect -60 785 180 790
rect -60 220 -15 785
rect 2 220 180 785
rect -60 215 180 220
rect 200 216 465 790
rect 485 216 666 791
rect 686 786 1196 791
rect 686 216 945 786
rect 200 215 945 216
rect -60 211 945 215
rect 965 211 1143 786
rect 1163 211 1196 786
rect -60 -8 1196 211
rect -60 -10 365 -8
rect -60 -585 -20 -10
rect 1 -583 365 -10
rect 386 -10 1196 -8
rect 386 -583 566 -10
rect 1 -585 566 -583
rect 587 -585 766 -10
rect 787 -14 1196 -10
rect 787 -585 1145 -14
rect -60 -589 1145 -585
rect 1166 -589 1196 -14
rect -60 -619 1196 -589
rect -60 -625 1090 -619
rect -60 -660 25 -625
rect 55 -654 1090 -625
rect 1120 -654 1196 -619
rect 55 -660 1196 -654
rect -60 -684 1196 -660
<< labels >>
rlabel metal1 -60 80 -60 80 7 VN
rlabel poly -90 44 -90 44 3 Vcn
rlabel poly -90 142 -90 142 3 Vbn
rlabel poly -90 950 -90 950 7 V2
rlabel poly -90 1655 -90 1655 7 V1
rlabel poly -90 1720 -90 1720 7 Vcp
rlabel metal1 -58 2455 -58 2455 7 Vp
rlabel poly -90 2475 -90 2475 7 Vbp
rlabel poly 1255 905 1255 905 3 Vout
<< end >>
