magic
tech sky130A
timestamp 1695781062
<< nwell >>
rect -70 270 85 950
<< nmos >>
rect 0 -185 15 215
rect 0 -360 15 -260
rect 0 -520 15 -420
<< pmos >>
rect 0 830 15 930
rect 0 670 15 770
rect 0 476 15 575
rect 0 290 15 390
<< ndiff >>
rect -50 195 0 215
rect -50 -165 -35 195
rect -15 -165 0 195
rect -50 -185 0 -165
rect 15 195 65 215
rect 15 -165 30 195
rect 50 -165 65 195
rect 15 -185 65 -165
rect -50 -280 0 -260
rect -50 -340 -35 -280
rect -15 -340 0 -280
rect -50 -360 0 -340
rect 15 -280 65 -260
rect 15 -340 30 -280
rect 50 -340 65 -280
rect 15 -360 65 -340
rect -50 -440 0 -420
rect -50 -500 -35 -440
rect -15 -500 0 -440
rect -50 -520 0 -500
rect 15 -440 65 -420
rect 15 -500 30 -440
rect 50 -500 65 -440
rect 15 -520 65 -500
<< pdiff >>
rect -50 910 0 930
rect -50 850 -35 910
rect -15 850 0 910
rect -50 830 0 850
rect 15 910 65 930
rect 15 850 30 910
rect 50 850 65 910
rect 15 830 65 850
rect -50 750 0 770
rect -50 690 -35 750
rect -15 690 0 750
rect -50 670 0 690
rect 15 750 65 770
rect 15 690 30 750
rect 50 690 65 750
rect 15 670 65 690
rect -50 555 0 575
rect -50 495 -35 555
rect -15 495 0 555
rect -50 476 0 495
rect 15 555 65 575
rect 15 495 30 555
rect 50 495 65 555
rect 15 476 65 495
rect -50 370 0 390
rect -50 310 -35 370
rect -15 310 0 370
rect -50 290 0 310
rect 15 370 65 390
rect 15 310 30 370
rect 50 310 65 370
rect 15 290 65 310
<< ndiffc >>
rect -35 -165 -15 195
rect 30 -165 50 195
rect -35 -340 -15 -280
rect 30 -340 50 -280
rect -35 -500 -15 -440
rect 30 -500 50 -440
<< pdiffc >>
rect -35 850 -15 910
rect 30 850 50 910
rect -35 690 -15 750
rect 30 690 50 750
rect -35 495 -15 555
rect 30 495 50 555
rect -35 310 -15 370
rect 30 310 50 370
<< poly >>
rect 0 930 15 945
rect 0 821 15 830
rect 0 820 80 821
rect 0 810 130 820
rect 0 806 80 810
rect 65 790 80 806
rect 100 804 130 810
rect 100 790 105 804
rect 0 770 15 785
rect 65 780 105 790
rect 0 655 15 670
rect -25 645 15 655
rect -25 625 -15 645
rect 5 625 15 645
rect -25 615 15 625
rect 0 575 15 588
rect -75 452 -41 460
rect -75 445 -66 452
rect -155 435 -66 445
rect -49 435 -41 452
rect -155 430 -41 435
rect -75 427 -41 430
rect 0 390 15 476
rect -65 266 -31 273
rect -65 255 -56 266
rect -135 249 -56 255
rect -39 249 -31 266
rect -135 240 -31 249
rect 0 215 15 290
rect 0 -200 15 -185
rect -115 -210 -78 -200
rect -115 -230 -105 -210
rect -86 -224 -78 -210
rect -86 -225 -55 -224
rect -86 -230 130 -225
rect -115 -240 130 -230
rect 0 -260 15 -240
rect 0 -374 15 -360
rect 65 -380 105 -370
rect 65 -395 75 -380
rect 0 -400 75 -395
rect 95 -400 105 -380
rect 0 -410 105 -400
rect 0 -420 15 -410
rect 0 -535 15 -520
<< polycont >>
rect 80 790 100 810
rect -15 625 5 645
rect -66 435 -49 452
rect -56 249 -39 266
rect -105 -230 -86 -210
rect 75 -400 95 -380
<< locali >>
rect -40 910 -10 920
rect -40 860 -35 910
rect -115 850 -35 860
rect -15 850 -10 910
rect -115 840 -10 850
rect 25 910 55 920
rect 25 850 30 910
rect 50 850 55 910
rect 25 840 55 850
rect -115 635 -95 840
rect 65 820 85 821
rect 65 810 105 820
rect 65 790 80 810
rect 100 790 105 810
rect 65 780 105 790
rect -40 750 -10 760
rect -40 690 -35 750
rect -15 690 -10 750
rect -40 680 -10 690
rect 25 750 55 760
rect 25 690 30 750
rect 50 690 55 750
rect 25 680 55 690
rect -25 645 15 655
rect -25 635 -15 645
rect -115 625 -15 635
rect 5 635 15 645
rect 5 625 55 635
rect -115 615 55 625
rect -115 -200 -95 615
rect 35 565 55 615
rect -40 555 -10 565
rect -40 495 -35 555
rect -15 495 -10 555
rect -40 485 -10 495
rect 25 555 55 565
rect 25 495 30 555
rect 50 495 55 555
rect 25 485 55 495
rect -40 462 -15 485
rect -58 460 -15 462
rect -75 452 -15 460
rect -75 435 -66 452
rect -49 445 -15 452
rect -49 435 -41 445
rect -75 427 -41 435
rect 85 425 105 780
rect 35 405 105 425
rect 35 380 55 405
rect -40 370 -10 380
rect -40 318 -35 370
rect -42 310 -35 318
rect -15 310 -10 370
rect -42 307 -10 310
rect -48 300 -10 307
rect 25 370 55 380
rect 25 310 30 370
rect 50 310 55 370
rect 25 300 55 310
rect -48 273 -25 300
rect -65 270 -25 273
rect -65 266 -31 270
rect -65 249 -56 266
rect -39 249 -31 266
rect -65 240 -31 249
rect -40 195 -10 205
rect -40 -165 -35 195
rect -15 -165 -10 195
rect -40 -175 -10 -165
rect 25 195 55 205
rect 25 -165 30 195
rect 50 -165 55 195
rect 25 -175 55 -165
rect -115 -210 -78 -200
rect -115 -230 -105 -210
rect -86 -230 -78 -210
rect -115 -240 -78 -230
rect -115 -540 -95 -240
rect -40 -270 -20 -175
rect 85 -270 105 405
rect -40 -280 -10 -270
rect -40 -340 -35 -280
rect -15 -340 -10 -280
rect -40 -350 -10 -340
rect 25 -280 105 -270
rect 25 -340 30 -280
rect 50 -290 105 -280
rect 50 -340 55 -290
rect 25 -350 55 -340
rect -40 -430 -20 -350
rect 85 -370 105 -290
rect 65 -380 105 -370
rect 65 -400 75 -380
rect 95 -400 105 -380
rect 65 -410 105 -400
rect -40 -440 -10 -430
rect -40 -500 -35 -440
rect -15 -500 -10 -440
rect -40 -510 -10 -500
rect 25 -440 55 -430
rect 25 -500 30 -440
rect 50 -500 55 -440
rect 25 -510 55 -500
rect 25 -540 45 -510
rect -115 -560 45 -540
<< end >>
