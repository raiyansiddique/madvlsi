magic
tech sky130A
timestamp 1695791791
<< nwell >>
rect -160 330 364 1010
<< nmos >>
rect 0 -185 15 215
rect 230 -10 245 90
rect 230 -160 245 -60
rect 0 -360 15 -260
rect 230 -380 245 -280
rect 0 -520 15 -420
rect 230 -540 245 -440
<< pmos >>
rect 0 890 15 990
rect 0 730 15 830
rect 230 735 245 835
rect 0 536 15 635
rect 230 535 245 635
rect 0 350 15 450
rect 230 350 245 450
<< ndiff >>
rect -50 195 0 215
rect -50 -165 -35 195
rect -15 -165 0 195
rect -50 -185 0 -165
rect 15 195 65 215
rect 15 -165 30 195
rect 50 -165 65 195
rect 180 70 230 90
rect 180 10 195 70
rect 215 10 230 70
rect 180 -10 230 10
rect 245 70 295 90
rect 245 10 260 70
rect 280 10 295 70
rect 245 -10 295 10
rect 180 -80 230 -60
rect 180 -140 195 -80
rect 215 -140 230 -80
rect 180 -160 230 -140
rect 245 -80 295 -60
rect 245 -140 260 -80
rect 280 -140 295 -80
rect 245 -160 295 -140
rect 15 -185 65 -165
rect -50 -280 0 -260
rect -50 -340 -35 -280
rect -15 -340 0 -280
rect -50 -360 0 -340
rect 15 -280 65 -260
rect 15 -340 30 -280
rect 50 -340 65 -280
rect 15 -360 65 -340
rect 180 -300 230 -280
rect 180 -360 195 -300
rect 215 -360 230 -300
rect 180 -380 230 -360
rect 245 -300 295 -280
rect 245 -360 260 -300
rect 280 -360 295 -300
rect 245 -380 295 -360
rect -50 -440 0 -420
rect -50 -500 -35 -440
rect -15 -500 0 -440
rect -50 -520 0 -500
rect 15 -440 65 -420
rect 15 -500 30 -440
rect 50 -500 65 -440
rect 15 -520 65 -500
rect 180 -460 230 -440
rect 180 -520 195 -460
rect 215 -520 230 -460
rect 180 -540 230 -520
rect 245 -460 295 -440
rect 245 -520 260 -460
rect 280 -520 295 -460
rect 245 -540 295 -520
<< pdiff >>
rect -50 970 0 990
rect -50 910 -35 970
rect -15 910 0 970
rect -50 890 0 910
rect 15 970 65 990
rect 15 910 30 970
rect 50 910 65 970
rect 15 890 65 910
rect -50 810 0 830
rect -50 750 -35 810
rect -15 750 0 810
rect -50 730 0 750
rect 15 810 65 830
rect 15 750 30 810
rect 50 750 65 810
rect 15 730 65 750
rect 180 815 230 835
rect 180 755 195 815
rect 215 755 230 815
rect 180 735 230 755
rect 245 815 295 835
rect 245 755 260 815
rect 280 755 295 815
rect 245 735 295 755
rect -50 615 0 635
rect -50 555 -35 615
rect -15 555 0 615
rect -50 536 0 555
rect 15 615 65 635
rect 15 555 30 615
rect 50 555 65 615
rect 15 536 65 555
rect 180 615 230 635
rect 180 555 195 615
rect 215 555 230 615
rect 180 535 230 555
rect 245 615 295 635
rect 245 555 260 615
rect 280 555 295 615
rect 245 535 295 555
rect -50 430 0 450
rect -50 370 -35 430
rect -15 370 0 430
rect -50 350 0 370
rect 15 430 65 450
rect 15 370 30 430
rect 50 370 65 430
rect 15 350 65 370
rect 180 430 230 450
rect 180 370 195 430
rect 215 370 230 430
rect 180 350 230 370
rect 245 430 295 450
rect 245 370 260 430
rect 280 370 295 430
rect 245 350 295 370
<< ndiffc >>
rect -35 -165 -15 195
rect 30 -165 50 195
rect 195 10 215 70
rect 260 10 280 70
rect 195 -140 215 -80
rect 260 -140 280 -80
rect -35 -340 -15 -280
rect 30 -340 50 -280
rect 195 -360 215 -300
rect 260 -360 280 -300
rect -35 -500 -15 -440
rect 30 -500 50 -440
rect 195 -520 215 -460
rect 260 -520 280 -460
<< pdiffc >>
rect -35 910 -15 970
rect 30 910 50 970
rect -35 750 -15 810
rect 30 750 50 810
rect 195 755 215 815
rect 260 755 280 815
rect -35 555 -15 615
rect 30 555 50 615
rect 195 555 215 615
rect 260 555 280 615
rect -35 370 -15 430
rect 30 370 50 430
rect 195 370 215 430
rect 260 370 280 430
<< psubdiff >>
rect 155 190 205 213
rect 155 140 173 190
rect 190 140 205 190
rect 155 121 205 140
<< nsubdiff >>
rect 196 970 246 992
rect 196 915 212 970
rect 229 915 246 970
rect 196 892 246 915
<< psubdiffcont >>
rect 173 140 190 190
<< nsubdiffcont >>
rect 212 915 229 970
<< poly >>
rect 0 990 15 1005
rect 0 881 15 890
rect 0 880 80 881
rect 0 870 105 880
rect 0 866 80 870
rect 65 850 80 866
rect 100 850 105 870
rect 0 830 15 845
rect 65 840 105 850
rect 230 835 245 848
rect 0 715 15 730
rect -25 705 15 715
rect -25 685 -15 705
rect 5 685 15 705
rect 230 716 245 735
rect 230 715 295 716
rect 230 705 320 715
rect 230 701 290 705
rect -25 675 15 685
rect 123 685 163 696
rect 123 665 134 685
rect 153 680 163 685
rect 280 685 290 701
rect 310 685 320 705
rect 153 665 245 680
rect 280 675 320 685
rect 123 663 245 665
rect 123 656 163 663
rect 0 635 15 648
rect -75 512 -41 520
rect -75 505 -66 512
rect -155 495 -66 505
rect -49 495 -41 512
rect -155 490 -41 495
rect -75 487 -41 490
rect 0 450 15 536
rect 123 500 140 656
rect 230 635 245 663
rect 230 522 245 535
rect 320 500 370 505
rect 123 490 370 500
rect 123 485 335 490
rect -65 326 -31 333
rect -65 315 -56 326
rect -155 309 -56 315
rect -39 309 -31 326
rect -155 300 -31 309
rect 0 280 15 350
rect -15 274 25 280
rect -15 257 -5 274
rect 16 257 25 274
rect -15 250 25 257
rect 0 215 15 250
rect 123 0 140 485
rect 230 450 245 463
rect 230 280 245 350
rect 305 315 345 320
rect 305 314 370 315
rect 305 297 315 314
rect 334 300 370 314
rect 334 297 345 300
rect 305 290 345 297
rect 220 274 260 280
rect 220 257 229 274
rect 250 257 260 274
rect 220 250 260 257
rect 230 90 245 250
rect 123 -10 163 0
rect 123 -30 135 -10
rect 154 -30 163 -10
rect 123 -40 163 -30
rect 230 -60 245 -10
rect 230 -173 245 -160
rect 0 -200 15 -185
rect -115 -210 -78 -200
rect -115 -230 -105 -210
rect -86 -224 -78 -210
rect 162 -205 202 -195
rect 162 -220 170 -205
rect -86 -225 -55 -224
rect 93 -225 170 -220
rect 190 -225 202 -205
rect 248 -205 285 -195
rect 248 -218 259 -205
rect -86 -230 202 -225
rect -115 -235 202 -230
rect 230 -225 259 -218
rect 276 -225 285 -205
rect 230 -235 285 -225
rect -115 -240 109 -235
rect 0 -260 15 -240
rect 230 -280 245 -235
rect 0 -374 15 -360
rect 65 -380 105 -370
rect 65 -395 75 -380
rect 0 -400 75 -395
rect 95 -400 105 -380
rect 230 -393 245 -380
rect 0 -410 105 -400
rect 0 -420 15 -410
rect 293 -417 330 -398
rect 230 -432 330 -417
rect 230 -440 245 -432
rect 0 -535 15 -520
rect 230 -557 245 -540
<< polycont >>
rect 80 850 100 870
rect -15 685 5 705
rect 134 665 153 685
rect 290 685 310 705
rect -66 495 -49 512
rect -56 309 -39 326
rect -5 257 16 274
rect 315 297 334 314
rect 229 257 250 274
rect 135 -30 154 -10
rect -105 -230 -86 -210
rect 170 -225 190 -205
rect 259 -225 276 -205
rect 75 -400 95 -380
<< locali >>
rect -40 970 -10 980
rect -40 920 -35 970
rect -115 910 -35 920
rect -15 910 -10 970
rect -115 900 -10 910
rect 25 970 55 980
rect 25 910 30 970
rect 50 910 55 970
rect 25 900 55 910
rect 205 970 235 980
rect 205 915 212 970
rect 229 915 235 970
rect 205 903 235 915
rect -115 695 -95 900
rect 65 880 85 881
rect 65 870 105 880
rect 65 850 80 870
rect 100 850 105 870
rect 65 840 105 850
rect 85 820 105 840
rect -40 810 -10 820
rect -40 750 -35 810
rect -15 750 -10 810
rect -40 740 -10 750
rect 25 810 105 820
rect 25 750 30 810
rect 50 800 105 810
rect 50 750 55 800
rect 25 740 55 750
rect -25 705 15 715
rect -25 695 -15 705
rect -115 685 -15 695
rect 5 695 15 705
rect 5 685 55 695
rect -115 675 55 685
rect -115 -200 -95 675
rect 35 625 55 675
rect -40 615 -10 625
rect -40 555 -35 615
rect -15 555 -10 615
rect -40 545 -10 555
rect 25 615 55 625
rect 25 555 30 615
rect 50 555 55 615
rect 25 545 55 555
rect -40 522 -15 545
rect -58 520 -15 522
rect -75 512 -15 520
rect -75 495 -66 512
rect -49 505 -15 512
rect -49 495 -41 505
rect -75 487 -41 495
rect 85 485 105 800
rect 123 865 275 885
rect 123 696 140 865
rect 255 825 275 865
rect 190 815 220 825
rect 190 755 195 815
rect 215 755 220 815
rect 190 745 220 755
rect 255 815 285 825
rect 255 755 260 815
rect 280 755 285 815
rect 255 745 285 755
rect 123 685 163 696
rect 123 665 134 685
rect 153 665 163 685
rect 123 656 163 665
rect 190 625 209 745
rect 280 705 330 715
rect 280 685 290 705
rect 310 685 330 705
rect 280 675 330 685
rect 190 615 220 625
rect 190 555 195 615
rect 215 555 220 615
rect 190 545 220 555
rect 255 615 285 625
rect 255 555 260 615
rect 280 565 285 615
rect 310 565 330 675
rect 280 555 330 565
rect 255 545 330 555
rect 35 465 105 485
rect 35 440 55 465
rect -40 430 -10 440
rect -40 378 -35 430
rect -42 370 -35 378
rect -15 370 -10 430
rect -42 367 -10 370
rect -48 360 -10 367
rect 25 430 55 440
rect 25 370 30 430
rect 50 370 55 430
rect 25 360 55 370
rect -48 333 -25 360
rect -65 330 -25 333
rect -65 326 -31 330
rect -65 309 -56 326
rect -39 309 -31 326
rect -65 300 -31 309
rect -15 274 25 280
rect -15 257 -5 274
rect 16 257 25 274
rect -15 250 25 257
rect -40 195 -10 205
rect -40 -165 -35 195
rect -15 -165 -10 195
rect -40 -175 -10 -165
rect 25 195 55 205
rect 25 -165 30 195
rect 50 -165 55 195
rect 25 -175 55 -165
rect 85 80 105 465
rect 191 440 210 545
rect 190 430 220 440
rect 190 370 195 430
rect 215 370 220 430
rect 190 360 220 370
rect 255 430 285 440
rect 255 370 260 430
rect 280 370 285 430
rect 255 360 285 370
rect 310 320 330 545
rect 305 314 345 320
rect 305 297 315 314
rect 334 297 345 314
rect 305 290 345 297
rect 220 274 260 280
rect 220 257 229 274
rect 250 257 260 274
rect 220 250 260 257
rect 165 190 195 200
rect 165 140 173 190
rect 190 140 195 190
rect 165 130 195 140
rect 310 80 330 290
rect 85 70 220 80
rect 85 60 195 70
rect -115 -210 -78 -200
rect -115 -230 -105 -210
rect -86 -230 -78 -210
rect -115 -240 -78 -230
rect -115 -540 -95 -240
rect -40 -270 -20 -175
rect 85 -270 105 60
rect 190 10 195 60
rect 215 10 220 70
rect 190 0 220 10
rect 255 70 330 80
rect 255 10 260 70
rect 280 60 330 70
rect 280 10 285 60
rect 255 0 285 10
rect -40 -280 -10 -270
rect -40 -340 -35 -280
rect -15 -340 -10 -280
rect -40 -350 -10 -340
rect 25 -280 105 -270
rect 123 -10 163 0
rect 123 -30 135 -10
rect 154 -30 163 -10
rect 123 -40 163 -30
rect 123 -252 143 -40
rect 190 -80 220 -70
rect 190 -132 195 -80
rect 185 -140 195 -132
rect 215 -140 220 -80
rect 185 -150 220 -140
rect 255 -80 285 -70
rect 255 -140 260 -80
rect 280 -140 285 -80
rect 255 -150 285 -140
rect 185 -195 202 -150
rect 265 -195 285 -150
rect 162 -205 202 -195
rect 162 -225 170 -205
rect 190 -225 202 -205
rect 162 -235 202 -225
rect 248 -205 285 -195
rect 248 -225 259 -205
rect 276 -225 285 -205
rect 248 -235 285 -225
rect 260 -252 280 -235
rect 123 -266 280 -252
rect 123 -270 271 -266
rect 123 -272 170 -270
rect 25 -340 30 -280
rect 50 -290 105 -280
rect 50 -340 55 -290
rect 25 -350 55 -340
rect -40 -430 -20 -350
rect 85 -370 105 -290
rect 65 -380 105 -370
rect 65 -400 75 -380
rect 95 -400 105 -380
rect 65 -410 105 -400
rect -40 -440 -10 -430
rect -40 -500 -35 -440
rect -15 -500 -10 -440
rect -40 -510 -10 -500
rect 25 -440 55 -430
rect 25 -500 30 -440
rect 50 -500 55 -440
rect 150 -455 170 -272
rect 310 -290 330 60
rect 190 -300 220 -290
rect 190 -360 195 -300
rect 215 -360 220 -300
rect 190 -370 220 -360
rect 255 -300 330 -290
rect 255 -360 260 -300
rect 280 -310 330 -300
rect 280 -360 285 -310
rect 255 -370 285 -360
rect 310 -398 330 -310
rect 293 -432 330 -398
rect 190 -455 220 -450
rect 150 -460 220 -455
rect 150 -474 195 -460
rect 25 -510 55 -500
rect 25 -540 45 -510
rect 190 -520 195 -474
rect 215 -520 220 -460
rect 190 -530 220 -520
rect 255 -460 285 -450
rect 255 -520 260 -460
rect 280 -520 285 -460
rect 255 -530 285 -520
rect -115 -560 45 -540
<< viali >>
rect 30 910 50 970
rect 212 915 229 970
rect -35 750 -15 810
rect -5 257 16 274
rect 30 -165 50 195
rect 260 370 280 430
rect 229 257 250 274
rect 173 140 190 190
rect 195 -360 215 -300
rect 260 -520 280 -460
<< metal1 >>
rect -145 970 355 1005
rect -145 910 30 970
rect 50 915 212 970
rect 229 915 355 970
rect 50 910 355 915
rect -145 810 355 910
rect -145 750 -35 810
rect -15 750 355 810
rect -145 430 355 750
rect -145 370 260 430
rect 280 370 355 430
rect -145 335 355 370
rect -145 274 350 280
rect -145 257 -5 274
rect 16 257 229 274
rect 250 257 350 274
rect -145 250 350 257
rect -145 195 350 220
rect -145 -165 30 195
rect 50 190 350 195
rect 50 140 173 190
rect 190 140 350 190
rect 50 -165 350 140
rect -145 -300 350 -165
rect -145 -360 195 -300
rect 215 -360 350 -300
rect -145 -460 350 -360
rect -145 -520 260 -460
rect 280 -520 350 -460
rect -145 -565 350 -520
<< labels >>
rlabel metal1 -145 640 -145 640 7 VP
port 2 w
rlabel metal1 -145 160 -145 160 7 VN
port 5 w
rlabel metal1 -145 265 -145 265 7 CLK
port 4 w
rlabel poly -155 308 -155 308 7 D_bar
port 3 w
rlabel poly -155 498 -155 498 7 D
port 1 w
rlabel poly 370 497 370 497 3 Q
port 7 e
rlabel poly 370 308 370 308 3 Q_bar
port 6 e
<< end >>
