* SPICE3 file created from buffer.ext - technology: sky130A

.subckt inverter A Y VP VN
X0 Y A VN VN sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.15
.ends

.subckt buffer
Xinverter_0 inverter_0/A inverter_1/A VN VP inverter
Xinverter_1 inverter_1/A Y VN VP inverter
.ends

