magic
tech sky130A
timestamp 1694659262
<< nwell >>
rect -75 150 200 300
<< nmos >>
rect 50 0 65 100
rect 115 0 130 100
<< pmos >>
rect 50 170 65 270
rect 115 170 130 270
<< ndiff >>
rect 0 85 50 100
rect 0 15 15 85
rect 35 15 50 85
rect 0 0 50 15
rect 65 0 115 100
rect 130 85 180 100
rect 130 15 145 85
rect 165 15 180 85
rect 130 0 180 15
<< pdiff >>
rect 0 255 50 270
rect 0 185 15 255
rect 35 185 50 255
rect 0 170 50 185
rect 65 255 115 270
rect 65 186 80 255
rect 100 186 115 255
rect 65 170 115 186
rect 130 255 180 270
rect 130 185 145 255
rect 165 185 180 255
rect 130 170 180 185
<< ndiffc >>
rect 15 15 35 85
rect 145 15 165 85
<< pdiffc >>
rect 15 185 35 255
rect 80 186 100 255
rect 145 185 165 255
<< psubdiff >>
rect -50 85 0 100
rect -50 15 -30 85
rect -10 15 0 85
rect -50 0 0 15
<< nsubdiff >>
rect -50 255 0 270
rect -50 185 -30 255
rect -10 185 0 255
rect -50 170 0 185
<< psubdiffcont >>
rect -30 15 -10 85
<< nsubdiffcont >>
rect -30 185 -10 255
<< poly >>
rect 50 270 65 293
rect 115 270 130 295
rect 50 100 65 170
rect 115 100 130 170
rect 50 -20 65 0
rect 25 -30 65 -20
rect 25 -50 35 -30
rect 55 -50 65 -30
rect 25 -60 65 -50
rect 115 -60 130 0
rect 90 -70 130 -60
rect 90 -90 100 -70
rect 120 -90 130 -70
rect 90 -100 130 -90
<< polycont >>
rect 35 -50 55 -30
rect 100 -90 120 -70
<< locali >>
rect -40 255 45 265
rect -40 185 -30 255
rect -10 185 15 255
rect 35 185 45 255
rect -40 175 45 185
rect 70 255 110 265
rect 70 186 80 255
rect 100 186 110 255
rect 70 175 110 186
rect 135 255 175 265
rect 135 185 145 255
rect 165 185 175 255
rect 135 175 175 185
rect 90 155 110 175
rect 90 135 200 155
rect 145 95 165 135
rect -40 85 45 95
rect -40 15 -30 85
rect -10 15 15 85
rect 35 15 45 85
rect -40 5 45 15
rect 135 85 175 95
rect 135 15 145 85
rect 165 15 175 85
rect 135 5 175 15
rect -75 -30 65 -20
rect -75 -40 35 -30
rect 25 -50 35 -40
rect 55 -50 65 -30
rect 25 -60 65 -50
rect 90 -70 130 -60
rect 90 -80 100 -70
rect -75 -90 100 -80
rect 120 -90 130 -70
rect -75 -100 130 -90
<< viali >>
rect -30 185 -10 255
rect 15 185 35 255
rect 145 185 165 255
rect -30 15 -10 85
rect 15 15 35 85
<< metal1 >>
rect -75 255 200 265
rect -75 185 -30 255
rect -10 185 15 255
rect 35 185 145 255
rect 165 185 200 255
rect -75 175 200 185
rect -75 85 200 95
rect -75 15 -30 85
rect -10 15 15 85
rect 35 15 200 85
rect -75 5 200 15
<< labels >>
rlabel metal1 -75 220 -75 220 7 VP
port 1 w
rlabel metal1 -75 50 -75 50 7 VN
port 2 w
rlabel locali -75 -30 -75 -30 7 A
port 3 w
rlabel locali -75 -90 -75 -90 7 B
port 4 w
rlabel locali 200 145 200 145 3 Y
port 5 e
<< end >>
