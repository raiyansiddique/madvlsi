magic
tech sky130A
timestamp 1697333037
<< error_p >>
rect 194 -4 195 12
rect 194 -21 195 -5
rect 606 -599 607 1
<< nmos >>
rect 0 -600 50 0
rect 100 -600 150 0
rect 200 -600 250 0
rect 381 -599 431 1
rect 481 -599 531 1
rect 656 -599 706 1
rect 756 -599 806 1
rect 856 -599 906 1
<< ndiff >>
rect -50 -10 0 0
rect -50 -585 -35 -10
rect -15 -585 0 -10
rect -50 -600 0 -585
rect 50 -10 100 0
rect 50 -585 65 -10
rect 85 -585 100 -10
rect 50 -600 100 -585
rect 150 -10 200 0
rect 150 -585 165 -10
rect 185 -585 200 -10
rect 150 -600 200 -585
rect 250 -10 300 0
rect 250 -585 265 -10
rect 285 -585 300 -10
rect 250 -600 300 -585
rect 331 -9 381 1
rect 331 -584 346 -9
rect 366 -584 381 -9
rect 331 -599 381 -584
rect 431 -9 481 1
rect 431 -584 446 -9
rect 466 -584 481 -9
rect 431 -599 481 -584
rect 531 -9 580 1
rect 531 -584 546 -9
rect 566 -584 580 -9
rect 531 -599 580 -584
rect 606 -9 656 1
rect 606 -584 621 -9
rect 641 -584 656 -9
rect 606 -599 656 -584
rect 706 -9 756 1
rect 706 -584 721 -9
rect 741 -584 756 -9
rect 706 -599 756 -584
rect 806 -9 856 1
rect 806 -584 821 -9
rect 841 -584 856 -9
rect 806 -599 856 -584
rect 906 -9 956 1
rect 906 -584 921 -9
rect 940 -584 956 -9
rect 906 -599 956 -584
<< ndiffc >>
rect -35 -585 -15 -10
rect 65 -585 85 -10
rect 165 -585 185 -10
rect 265 -585 285 -10
rect 346 -584 366 -9
rect 446 -584 466 -9
rect 546 -584 566 -9
rect 621 -584 641 -9
rect 721 -584 741 -9
rect 821 -584 841 -9
rect 921 -584 940 -9
<< poly >>
rect 0 55 50 65
rect 0 20 10 55
rect 40 20 50 55
rect 0 0 50 20
rect 100 0 150 13
rect 200 0 250 13
rect 381 1 431 14
rect 481 1 531 14
rect 656 1 706 14
rect 756 1 806 14
rect 856 1 906 14
rect 0 -615 50 -600
rect 100 -615 150 -600
rect 200 -615 250 -600
rect 381 -614 431 -599
rect 481 -614 531 -599
rect 656 -614 706 -599
rect 756 -614 806 -599
rect 856 -615 906 -599
<< polycont >>
rect 10 20 40 55
<< locali >>
rect 0 55 50 65
rect 0 20 10 55
rect 40 20 50 55
rect 0 13 50 20
rect 155 30 475 55
rect 155 0 195 30
rect 154 -4 195 0
rect 154 -5 194 -4
rect -45 -10 -5 -5
rect -45 -585 -35 -10
rect -15 -585 -5 -10
rect -45 -595 -5 -585
rect 55 -10 95 -5
rect 55 -585 65 -10
rect 85 -585 95 -10
rect 154 -10 195 -5
rect 154 -27 165 -10
rect 55 -591 95 -585
rect 155 -585 165 -27
rect 185 -585 195 -10
rect 55 -625 96 -591
rect 155 -595 195 -585
rect 255 -10 295 -5
rect 255 -585 265 -10
rect 285 -585 295 -10
rect 255 -625 295 -585
rect 55 -652 295 -625
rect 336 -9 376 1
rect 336 -584 346 -9
rect 366 -584 376 -9
rect 435 -4 475 30
rect 435 -9 476 -4
rect 435 -10 446 -9
rect 336 -594 376 -584
rect 436 -584 446 -10
rect 466 -584 476 -9
rect 436 -594 476 -584
rect 536 -9 576 -4
rect 536 -584 546 -9
rect 566 -584 576 -9
rect 536 -594 576 -584
rect 611 -9 651 -4
rect 611 -584 621 -9
rect 641 -584 651 -9
rect 611 -594 651 -584
rect 711 -9 751 -4
rect 711 -584 721 -9
rect 741 -584 751 -9
rect 711 -594 751 -584
rect 811 -9 851 -4
rect 811 -584 821 -9
rect 841 -584 851 -9
rect 811 -594 851 -584
rect 911 -9 951 -4
rect 911 -584 921 -9
rect 940 -584 951 -9
rect 911 -594 951 -584
rect 336 -625 375 -594
rect 436 -599 475 -594
rect 536 -625 575 -594
rect 336 -650 575 -625
rect 336 -651 475 -650
<< end >>
