** sch_path: /home/madvlsi/madvlsi/mp1/cmos_inverter/buffer.sch
**.subckt buffer A VP VN Y
*.ipin A
*.iopin VP
*.iopin VN
*.opin Y
X1 A VN VP net1 inverter
X2 net1 VN VP Y inverter
**.ends

* expanding   symbol:  /home/madvlsi/madvlsi/mp1/cmos_inverter/inverter.sym # of pins=4
** sym_path: /home/madvlsi/madvlsi/mp1/cmos_inverter/inverter.sym
** sch_path: /home/madvlsi/madvlsi/mp1/cmos_inverter/inverter.sch
.subckt inverter A VN VP Y
*.ipin A
*.iopin VP
*.iopin VN
*.opin Y
XM1 Y A VN VN sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Y A VP VP sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
