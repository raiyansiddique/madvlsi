magic
tech sky130A
timestamp 1697429042
<< nwell >>
rect -277 1021 1788 2556
<< nmos >>
rect 0 150 50 750
rect 100 150 150 750
rect 200 150 250 750
rect 300 150 350 750
rect 400 150 450 750
rect 500 150 550 750
rect 600 150 650 750
rect 700 150 750 750
rect 800 150 850 750
rect 900 150 950 750
rect 1000 150 1050 750
rect 1100 150 1150 750
rect 1200 150 1250 750
rect 1300 150 1350 750
rect 1400 150 1450 750
rect 1500 150 1550 750
rect 0 -600 50 0
rect 100 -600 150 0
rect 200 -600 250 0
rect 300 -600 350 0
rect 400 -600 450 0
rect 500 -600 550 0
rect 600 -600 650 0
rect 700 -600 750 0
rect 800 -600 850 0
rect 900 -600 950 0
rect 1000 -600 1050 0
rect 1100 -600 1150 0
rect 1200 -600 1250 0
rect 1300 -600 1350 0
rect 1400 -600 1450 0
rect 1500 -600 1550 0
<< pmos >>
rect 0 1875 50 2475
rect 100 1875 150 2475
rect 200 1875 250 2475
rect 300 1875 350 2475
rect 400 1875 450 2475
rect 500 1875 550 2475
rect 600 1875 650 2475
rect 700 1875 750 2475
rect 800 1875 850 2475
rect 900 1875 950 2475
rect 1000 1875 1050 2475
rect 1100 1875 1150 2475
rect 1200 1875 1250 2475
rect 1300 1875 1350 2475
rect 1400 1875 1450 2475
rect 1500 1875 1550 2475
rect 0 1125 50 1725
rect 100 1125 150 1725
rect 200 1125 250 1725
rect 300 1125 350 1725
rect 400 1125 450 1725
rect 500 1125 550 1725
rect 600 1125 650 1725
rect 700 1125 750 1725
rect 800 1125 850 1725
rect 900 1125 950 1725
rect 1000 1125 1050 1725
rect 1100 1125 1150 1725
rect 1200 1125 1250 1725
rect 1300 1125 1350 1725
rect 1400 1125 1450 1725
rect 1500 1125 1550 1725
<< ndiff >>
rect -50 735 0 750
rect -50 165 -35 735
rect -15 165 0 735
rect -50 150 0 165
rect 50 735 100 750
rect 50 165 65 735
rect 85 165 100 735
rect 50 150 100 165
rect 150 735 200 750
rect 150 165 165 735
rect 185 165 200 735
rect 150 150 200 165
rect 250 735 300 750
rect 250 165 265 735
rect 285 165 300 735
rect 250 150 300 165
rect 350 735 400 750
rect 350 165 365 735
rect 385 165 400 735
rect 350 150 400 165
rect 450 735 500 750
rect 450 165 465 735
rect 485 165 500 735
rect 450 150 500 165
rect 550 735 600 750
rect 550 165 565 735
rect 585 165 600 735
rect 550 150 600 165
rect 650 735 700 750
rect 650 165 665 735
rect 685 165 700 735
rect 650 150 700 165
rect 750 735 800 750
rect 750 165 765 735
rect 785 165 800 735
rect 750 150 800 165
rect 850 735 900 750
rect 850 165 865 735
rect 885 165 900 735
rect 850 150 900 165
rect 950 735 1000 750
rect 950 165 965 735
rect 985 165 1000 735
rect 950 150 1000 165
rect 1050 735 1100 750
rect 1050 165 1065 735
rect 1085 165 1100 735
rect 1050 150 1100 165
rect 1150 735 1200 750
rect 1150 165 1165 735
rect 1185 165 1200 735
rect 1150 150 1200 165
rect 1250 735 1300 750
rect 1250 165 1265 735
rect 1285 165 1300 735
rect 1250 150 1300 165
rect 1350 735 1400 750
rect 1350 165 1365 735
rect 1385 165 1400 735
rect 1350 150 1400 165
rect 1450 735 1500 750
rect 1450 165 1465 735
rect 1485 165 1500 735
rect 1450 150 1500 165
rect 1550 735 1600 750
rect 1550 165 1565 735
rect 1585 165 1600 735
rect 1550 150 1600 165
rect -50 -15 0 0
rect -50 -585 -35 -15
rect -15 -585 0 -15
rect -50 -600 0 -585
rect 50 -15 100 0
rect 50 -585 65 -15
rect 85 -585 100 -15
rect 50 -600 100 -585
rect 150 -15 200 0
rect 150 -585 165 -15
rect 185 -585 200 -15
rect 150 -600 200 -585
rect 250 -15 300 0
rect 250 -585 265 -15
rect 285 -585 300 -15
rect 250 -600 300 -585
rect 350 -15 400 0
rect 350 -585 365 -15
rect 385 -585 400 -15
rect 350 -600 400 -585
rect 450 -15 500 0
rect 450 -585 465 -15
rect 485 -585 500 -15
rect 450 -600 500 -585
rect 550 -15 600 0
rect 550 -585 565 -15
rect 585 -585 600 -15
rect 550 -600 600 -585
rect 650 -15 700 0
rect 650 -585 665 -15
rect 685 -585 700 -15
rect 650 -600 700 -585
rect 750 -15 800 0
rect 750 -585 765 -15
rect 785 -585 800 -15
rect 750 -600 800 -585
rect 850 -15 900 0
rect 850 -585 865 -15
rect 885 -585 900 -15
rect 850 -600 900 -585
rect 950 -15 1000 0
rect 950 -585 965 -15
rect 985 -585 1000 -15
rect 950 -600 1000 -585
rect 1050 -15 1100 0
rect 1050 -585 1065 -15
rect 1085 -585 1100 -15
rect 1050 -600 1100 -585
rect 1150 -15 1200 0
rect 1150 -585 1165 -15
rect 1185 -585 1200 -15
rect 1150 -600 1200 -585
rect 1250 -15 1300 0
rect 1250 -585 1265 -15
rect 1285 -585 1300 -15
rect 1250 -600 1300 -585
rect 1350 -15 1400 0
rect 1350 -585 1365 -15
rect 1385 -585 1400 -15
rect 1350 -600 1400 -585
rect 1450 -15 1500 0
rect 1450 -585 1465 -15
rect 1485 -585 1500 -15
rect 1450 -600 1500 -585
rect 1550 -15 1600 0
rect 1550 -585 1565 -15
rect 1585 -585 1600 -15
rect 1550 -600 1600 -585
<< pdiff >>
rect -50 2460 0 2475
rect -50 1890 -35 2460
rect -15 1890 0 2460
rect -50 1875 0 1890
rect 50 2460 100 2475
rect 50 1890 65 2460
rect 85 1890 100 2460
rect 50 1875 100 1890
rect 150 2460 200 2475
rect 150 1890 165 2460
rect 185 1890 200 2460
rect 150 1875 200 1890
rect 250 2460 300 2475
rect 250 1890 265 2460
rect 285 1890 300 2460
rect 250 1875 300 1890
rect 350 2460 400 2475
rect 350 1890 365 2460
rect 385 1890 400 2460
rect 350 1875 400 1890
rect 450 2460 500 2475
rect 450 1890 465 2460
rect 485 1890 500 2460
rect 450 1875 500 1890
rect 550 2460 600 2475
rect 550 1890 565 2460
rect 585 1890 600 2460
rect 550 1875 600 1890
rect 650 2460 700 2475
rect 650 1890 665 2460
rect 685 1890 700 2460
rect 650 1875 700 1890
rect 750 2460 800 2475
rect 750 1890 765 2460
rect 785 1890 800 2460
rect 750 1875 800 1890
rect 850 2460 900 2475
rect 850 1890 865 2460
rect 885 1890 900 2460
rect 850 1875 900 1890
rect 950 2460 1000 2475
rect 950 1890 965 2460
rect 985 1890 1000 2460
rect 950 1875 1000 1890
rect 1050 2460 1100 2475
rect 1050 1890 1065 2460
rect 1085 1890 1100 2460
rect 1050 1875 1100 1890
rect 1150 2460 1200 2475
rect 1150 1890 1165 2460
rect 1185 1890 1200 2460
rect 1150 1875 1200 1890
rect 1250 2460 1300 2475
rect 1250 1890 1265 2460
rect 1285 1890 1300 2460
rect 1250 1875 1300 1890
rect 1350 2460 1400 2475
rect 1350 1890 1365 2460
rect 1385 1890 1400 2460
rect 1350 1875 1400 1890
rect 1450 2460 1500 2475
rect 1450 1890 1465 2460
rect 1485 1890 1500 2460
rect 1450 1875 1500 1890
rect 1550 2460 1600 2475
rect 1550 1890 1565 2460
rect 1585 1890 1600 2460
rect 1550 1875 1600 1890
rect -50 1710 0 1725
rect -50 1140 -35 1710
rect -15 1140 0 1710
rect -50 1125 0 1140
rect 50 1710 100 1725
rect 50 1140 65 1710
rect 85 1140 100 1710
rect 50 1125 100 1140
rect 150 1710 200 1725
rect 150 1140 165 1710
rect 185 1140 200 1710
rect 150 1125 200 1140
rect 250 1710 300 1725
rect 250 1140 265 1710
rect 285 1140 300 1710
rect 250 1125 300 1140
rect 350 1710 400 1725
rect 350 1140 365 1710
rect 385 1140 400 1710
rect 350 1125 400 1140
rect 450 1710 500 1725
rect 450 1140 465 1710
rect 485 1140 500 1710
rect 450 1125 500 1140
rect 550 1710 600 1725
rect 550 1140 565 1710
rect 585 1140 600 1710
rect 550 1125 600 1140
rect 650 1710 700 1725
rect 650 1140 665 1710
rect 685 1140 700 1710
rect 650 1125 700 1140
rect 750 1710 800 1725
rect 750 1140 765 1710
rect 785 1140 800 1710
rect 750 1125 800 1140
rect 850 1710 900 1725
rect 850 1140 865 1710
rect 885 1140 900 1710
rect 850 1125 900 1140
rect 950 1710 1000 1725
rect 950 1140 965 1710
rect 985 1140 1000 1710
rect 950 1125 1000 1140
rect 1050 1710 1100 1725
rect 1050 1140 1065 1710
rect 1085 1140 1100 1710
rect 1050 1125 1100 1140
rect 1150 1710 1200 1725
rect 1150 1140 1165 1710
rect 1185 1140 1200 1710
rect 1150 1125 1200 1140
rect 1250 1710 1300 1725
rect 1250 1140 1265 1710
rect 1285 1140 1300 1710
rect 1250 1125 1300 1140
rect 1350 1710 1400 1725
rect 1350 1140 1365 1710
rect 1385 1140 1400 1710
rect 1350 1125 1400 1140
rect 1450 1710 1500 1725
rect 1450 1140 1465 1710
rect 1485 1140 1500 1710
rect 1450 1125 1500 1140
rect 1550 1710 1600 1725
rect 1550 1140 1565 1710
rect 1585 1140 1600 1710
rect 1550 1125 1600 1140
<< ndiffc >>
rect -35 165 -15 735
rect 65 165 85 735
rect 165 165 185 735
rect 265 165 285 735
rect 365 165 385 735
rect 465 165 485 735
rect 565 165 585 735
rect 665 165 685 735
rect 765 165 785 735
rect 865 165 885 735
rect 965 165 985 735
rect 1065 165 1085 735
rect 1165 165 1185 735
rect 1265 165 1285 735
rect 1365 165 1385 735
rect 1465 165 1485 735
rect 1565 165 1585 735
rect -35 -585 -15 -15
rect 65 -585 85 -15
rect 165 -585 185 -15
rect 265 -585 285 -15
rect 365 -585 385 -15
rect 465 -585 485 -15
rect 565 -585 585 -15
rect 665 -585 685 -15
rect 765 -585 785 -15
rect 865 -585 885 -15
rect 965 -585 985 -15
rect 1065 -585 1085 -15
rect 1165 -585 1185 -15
rect 1265 -585 1285 -15
rect 1365 -585 1385 -15
rect 1465 -585 1485 -15
rect 1565 -585 1585 -15
<< pdiffc >>
rect -35 1890 -15 2460
rect 65 1890 85 2460
rect 165 1890 185 2460
rect 265 1890 285 2460
rect 365 1890 385 2460
rect 465 1890 485 2460
rect 565 1890 585 2460
rect 665 1890 685 2460
rect 765 1890 785 2460
rect 865 1890 885 2460
rect 965 1890 985 2460
rect 1065 1890 1085 2460
rect 1165 1890 1185 2460
rect 1265 1890 1285 2460
rect 1365 1890 1385 2460
rect 1465 1890 1485 2460
rect 1565 1890 1585 2460
rect -35 1140 -15 1710
rect 65 1140 85 1710
rect 165 1140 185 1710
rect 265 1140 285 1710
rect 365 1140 385 1710
rect 465 1140 485 1710
rect 565 1140 585 1710
rect 665 1140 685 1710
rect 765 1140 785 1710
rect 865 1140 885 1710
rect 965 1140 985 1710
rect 1065 1140 1085 1710
rect 1165 1140 1185 1710
rect 1265 1140 1285 1710
rect 1365 1140 1385 1710
rect 1465 1140 1485 1710
rect 1565 1140 1585 1710
<< psubdiff >>
rect -100 737 -50 750
rect -100 166 -90 737
rect -70 166 -50 737
rect -100 150 -50 166
rect 1600 735 1650 750
rect 1600 164 1620 735
rect 1640 164 1650 735
rect 1600 150 1650 164
rect -100 -15 -50 0
rect -100 -586 -90 -15
rect -70 -586 -50 -15
rect -100 -600 -50 -586
rect 1600 -14 1650 0
rect 1600 -585 1620 -14
rect 1640 -585 1650 -14
rect 1600 -600 1650 -585
<< nsubdiff >>
rect -100 2460 -50 2475
rect -100 1889 -90 2460
rect -70 1889 -50 2460
rect -100 1875 -50 1889
rect 1600 2461 1650 2475
rect 1600 1890 1620 2461
rect 1640 1890 1650 2461
rect 1600 1875 1650 1890
rect -100 1711 -50 1725
rect -100 1140 -90 1711
rect -70 1140 -50 1711
rect -100 1125 -50 1140
rect 1600 1709 1650 1725
rect 1600 1138 1620 1709
rect 1640 1138 1650 1709
rect 1600 1125 1650 1138
<< psubdiffcont >>
rect -90 166 -70 737
rect 1620 164 1640 735
rect -90 -586 -70 -15
rect 1620 -585 1640 -14
<< nsubdiffcont >>
rect -90 1889 -70 2460
rect 1620 1890 1640 2461
rect -90 1140 -70 1711
rect 1620 1138 1640 1709
<< poly >>
rect 1401 2591 2001 2630
rect 0 2520 50 2530
rect 0 2500 10 2520
rect 40 2500 50 2520
rect 1402 2517 1452 2591
rect 1300 2516 1452 2517
rect 0 2475 50 2500
rect 100 2490 1452 2516
rect 100 2475 150 2490
rect 200 2475 250 2490
rect 300 2475 350 2490
rect 400 2475 450 2490
rect 500 2475 550 2490
rect 600 2475 650 2490
rect 700 2475 750 2490
rect 800 2475 850 2490
rect 900 2475 950 2490
rect 1000 2475 1050 2490
rect 1100 2475 1150 2490
rect 1200 2475 1250 2490
rect 1300 2486 1452 2490
rect 1500 2520 1550 2529
rect 1500 2500 1510 2520
rect 1540 2500 1550 2520
rect 1300 2485 1450 2486
rect 1300 2475 1350 2485
rect 1400 2475 1450 2485
rect 1500 2475 1550 2500
rect 0 1725 50 1875
rect 100 1860 150 1875
rect 200 1860 250 1875
rect 300 1860 350 1875
rect 400 1860 450 1875
rect 500 1860 550 1875
rect 600 1860 650 1875
rect 700 1860 750 1875
rect 100 1775 150 1785
rect 800 1780 850 1875
rect 900 1860 950 1875
rect 1000 1860 1050 1875
rect 1100 1860 1150 1875
rect 1200 1860 1250 1875
rect 1300 1860 1350 1875
rect 1400 1860 1450 1875
rect 742 1778 850 1780
rect 100 1750 110 1775
rect 140 1750 150 1775
rect 100 1725 150 1750
rect 699 1770 850 1778
rect 699 1750 760 1770
rect 790 1750 850 1770
rect 699 1740 850 1750
rect 1400 1775 1450 1785
rect 1400 1750 1410 1775
rect 1440 1750 1450 1775
rect 200 1725 250 1740
rect 300 1725 350 1740
rect 400 1725 450 1740
rect 500 1725 550 1740
rect 600 1725 650 1740
rect 700 1725 750 1740
rect 800 1725 850 1740
rect 900 1725 950 1740
rect 1000 1725 1050 1740
rect 1100 1725 1150 1740
rect 1200 1725 1250 1740
rect 1300 1725 1350 1740
rect 1400 1725 1450 1750
rect 1500 1725 1550 1875
rect 0 1110 50 1125
rect 100 1110 150 1125
rect 200 1110 250 1125
rect 300 1110 350 1125
rect 400 1110 450 1125
rect 500 1110 550 1125
rect 600 1110 650 1125
rect 700 1110 750 1125
rect 800 1110 850 1125
rect 900 1110 950 1125
rect 1000 1110 1050 1125
rect 1100 1110 1150 1125
rect 1200 1110 1250 1125
rect 1300 1110 1350 1125
rect 1400 1110 1450 1125
rect 1500 1110 1550 1125
rect 101 990 148 1110
rect 210 1070 240 1110
rect 310 1070 340 1110
rect 410 1070 440 1110
rect 510 1070 540 1110
rect 610 1070 640 1110
rect 910 1070 940 1110
rect 1010 1070 1040 1110
rect 1110 1070 1140 1110
rect 1210 1070 1240 1110
rect 1310 1088 1340 1110
rect 1310 1079 1380 1088
rect 1310 1070 1350 1079
rect 200 1055 1350 1070
rect 1370 1055 1380 1079
rect 200 1045 1380 1055
rect 1415 990 1436 1110
rect 1775 990 1810 995
rect 101 987 1818 990
rect 101 971 1782 987
rect 1775 969 1782 971
rect 1801 971 1818 987
rect 1801 969 1810 971
rect 1775 959 1810 969
rect 1706 935 1753 948
rect -223 920 1724 935
rect -223 646 -207 920
rect 1706 915 1724 920
rect 1745 915 1753 935
rect 1706 907 1753 915
rect 100 869 1806 884
rect 100 765 127 869
rect 170 820 1350 830
rect 170 796 180 820
rect 200 805 1350 820
rect 200 796 240 805
rect 170 787 240 796
rect 210 765 240 787
rect 310 765 340 805
rect 410 765 440 805
rect 510 765 540 805
rect 610 765 640 805
rect 910 765 940 805
rect 1010 765 1040 805
rect 1110 765 1140 805
rect 1210 765 1240 805
rect 1310 765 1340 805
rect 1407 765 1445 869
rect 1743 868 1801 869
rect 0 750 50 765
rect 100 750 150 765
rect 200 750 250 765
rect 300 750 350 765
rect 400 750 450 765
rect 500 750 550 765
rect 600 750 650 765
rect 700 750 750 765
rect 800 750 850 765
rect 900 750 950 765
rect 1000 750 1050 765
rect 1100 750 1150 765
rect 1200 750 1250 765
rect 1300 750 1350 765
rect 1400 750 1450 765
rect 1500 750 1550 765
rect -223 635 -178 646
rect -223 616 -215 635
rect -186 616 -178 635
rect -223 608 -178 616
rect 0 0 50 150
rect 100 125 150 150
rect 200 135 250 150
rect 300 135 350 150
rect 400 135 450 150
rect 500 135 550 150
rect 600 135 650 150
rect 700 135 750 150
rect 800 135 850 150
rect 900 135 950 150
rect 1000 135 1050 150
rect 1100 135 1150 150
rect 1200 135 1250 150
rect 1300 135 1350 150
rect 100 100 110 125
rect 140 100 150 125
rect 100 90 150 100
rect 700 114 851 135
rect 1400 125 1450 150
rect 100 0 150 15
rect 200 0 250 15
rect 300 0 350 15
rect 400 0 450 15
rect 500 0 550 15
rect 600 0 650 15
rect 700 0 750 114
rect 1400 100 1410 125
rect 1440 100 1450 125
rect 1400 90 1450 100
rect 800 0 850 15
rect 900 0 950 15
rect 1000 0 1050 15
rect 1100 0 1150 15
rect 1200 0 1250 15
rect 1300 0 1350 15
rect 1400 0 1450 15
rect 1500 0 1550 150
rect 0 -625 50 -600
rect 100 -610 150 -600
rect 200 -610 250 -600
rect 100 -614 250 -610
rect 0 -645 10 -625
rect 40 -645 50 -625
rect 101 -615 250 -614
rect 300 -615 350 -600
rect 400 -615 450 -600
rect 500 -615 550 -600
rect 600 -615 650 -600
rect 700 -615 750 -600
rect 800 -615 850 -600
rect 900 -615 950 -600
rect 1000 -615 1050 -600
rect 1100 -615 1150 -600
rect 1200 -615 1250 -600
rect 1300 -615 1350 -600
rect 1400 -615 1450 -600
rect 101 -641 1450 -615
rect 1500 -625 1550 -600
rect 101 -642 250 -641
rect 0 -654 50 -645
rect 99 -682 128 -642
rect 1500 -645 1510 -625
rect 1540 -645 1550 -625
rect 1500 -655 1550 -645
rect -243 -708 128 -682
rect -243 -709 126 -708
<< polycont >>
rect 10 2500 40 2520
rect 1510 2500 1540 2520
rect 110 1750 140 1775
rect 760 1750 790 1770
rect 1410 1750 1440 1775
rect 1350 1055 1370 1079
rect 1782 969 1801 987
rect 1724 915 1745 935
rect 180 796 200 820
rect -215 616 -186 635
rect 110 100 140 125
rect 1410 100 1440 125
rect 10 -645 40 -625
rect 1510 -645 1540 -625
<< locali >>
rect -193 2563 92 2564
rect -193 2562 1480 2563
rect -195 2552 1480 2562
rect -195 2547 1481 2552
rect -195 2509 -175 2547
rect 69 2542 1481 2547
rect 0 2520 50 2530
rect -194 2484 -176 2509
rect 0 2500 10 2520
rect 40 2500 50 2520
rect 0 2490 50 2500
rect 69 2525 92 2542
rect -194 2362 -174 2484
rect -45 2470 -25 2473
rect -195 2251 -174 2362
rect -95 2460 -64 2470
rect -195 786 -175 2251
rect -95 1889 -90 2460
rect -70 1889 -64 2460
rect -95 1880 -64 1889
rect -45 2460 -5 2470
rect 69 2467 91 2525
rect 1455 2470 1481 2542
rect 1500 2520 1550 2529
rect 1500 2500 1510 2520
rect 1540 2500 1550 2520
rect 1500 2490 1550 2500
rect 69 2465 95 2467
rect -45 1890 -35 2460
rect -15 1890 -5 2460
rect -45 1880 -5 1890
rect 55 2460 95 2465
rect 55 1890 65 2460
rect 85 1890 95 2460
rect 55 1880 95 1890
rect 155 2461 195 2470
rect 155 1890 165 2461
rect 185 1890 195 2461
rect 155 1880 195 1890
rect 255 2460 295 2470
rect 255 1890 265 2460
rect 285 1890 295 2460
rect 255 1880 295 1890
rect 355 2460 395 2470
rect 355 1890 365 2460
rect 385 1890 395 2460
rect 355 1880 395 1890
rect 455 2460 495 2470
rect 455 1890 465 2460
rect 485 1890 495 2460
rect 455 1880 495 1890
rect 555 2460 595 2470
rect 555 1890 565 2460
rect 585 1890 595 2460
rect 555 1880 595 1890
rect 655 2460 695 2470
rect 655 1890 665 2460
rect 685 1890 695 2460
rect 655 1880 695 1890
rect 755 2460 795 2470
rect 755 1890 765 2460
rect 785 1890 795 2460
rect 755 1880 795 1890
rect 855 2460 895 2470
rect 855 1890 865 2460
rect 885 1890 895 2460
rect 855 1880 895 1890
rect 955 2460 995 2470
rect 955 1890 965 2460
rect 985 1890 995 2460
rect 955 1880 995 1890
rect 1055 2460 1095 2470
rect 1055 1890 1065 2460
rect 1085 1890 1095 2460
rect 1055 1880 1095 1890
rect 1155 2460 1195 2470
rect 1155 1890 1165 2460
rect 1185 1890 1195 2460
rect 1155 1880 1195 1890
rect 1255 2460 1295 2470
rect 1255 1890 1265 2460
rect 1285 1890 1295 2460
rect 1255 1880 1295 1890
rect 1355 2460 1395 2470
rect 1355 1890 1365 2460
rect 1385 2459 1395 2460
rect 1355 1889 1366 1890
rect 1386 1889 1395 2459
rect 1355 1880 1395 1889
rect 1455 2460 1495 2470
rect 1455 1890 1465 2460
rect 1485 1890 1495 2460
rect 1455 1880 1495 1890
rect 1555 2460 1595 2470
rect 1555 1890 1565 2460
rect 1585 1890 1595 2460
rect 1555 1880 1595 1890
rect 1614 2461 1645 2470
rect 1614 1890 1620 2461
rect 1640 1890 1645 2461
rect 1614 1880 1645 1890
rect -152 1830 -127 1833
rect 755 1830 775 1880
rect -152 1805 776 1830
rect 1685 1825 1756 1826
rect 1478 1824 1756 1825
rect 795 1806 1756 1824
rect 795 1805 1620 1806
rect 1685 1805 1756 1806
rect -152 828 -127 1805
rect 63 1775 150 1785
rect 795 1780 812 1805
rect 742 1778 812 1780
rect 63 1765 110 1775
rect 63 1720 83 1765
rect 100 1750 110 1765
rect 140 1750 150 1775
rect 699 1770 848 1778
rect 100 1740 150 1750
rect 167 1745 594 1765
rect 167 1720 190 1745
rect 370 1720 395 1745
rect 569 1720 594 1745
rect 699 1750 760 1770
rect 790 1750 848 1770
rect 1400 1775 1490 1785
rect 699 1742 848 1750
rect 955 1747 1382 1764
rect 750 1740 803 1742
rect 760 1720 777 1740
rect 955 1720 985 1747
rect 1159 1720 1190 1747
rect 1365 1724 1382 1747
rect 1400 1750 1410 1775
rect 1440 1765 1490 1775
rect 1440 1750 1450 1765
rect 1400 1740 1450 1750
rect 1365 1720 1385 1724
rect 1470 1720 1490 1765
rect -95 1711 -64 1720
rect -95 1139 -90 1711
rect -70 1139 -64 1711
rect -95 1130 -64 1139
rect -45 1710 -5 1720
rect -45 1140 -35 1710
rect -15 1140 -5 1710
rect -45 1130 -5 1140
rect 55 1710 95 1720
rect 55 1140 65 1710
rect 85 1140 95 1710
rect 55 1130 95 1140
rect 155 1710 195 1720
rect 155 1140 165 1710
rect 185 1140 195 1710
rect 155 1130 195 1140
rect 255 1710 295 1720
rect 255 1140 265 1710
rect 285 1140 295 1710
rect 255 1130 295 1140
rect 355 1710 395 1720
rect 355 1140 365 1710
rect 385 1140 395 1710
rect 355 1130 395 1140
rect 455 1710 495 1720
rect 455 1140 465 1710
rect 485 1140 495 1710
rect 455 1130 495 1140
rect 555 1710 595 1720
rect 555 1140 565 1710
rect 585 1140 595 1710
rect 555 1130 595 1140
rect 655 1710 695 1720
rect 655 1140 665 1710
rect 685 1709 695 1710
rect 655 1139 666 1140
rect 686 1139 695 1709
rect 655 1130 695 1139
rect 755 1710 795 1720
rect 755 1140 765 1710
rect 785 1140 795 1710
rect 755 1130 795 1140
rect 855 1710 895 1720
rect 855 1140 865 1710
rect 885 1709 895 1710
rect 855 1139 866 1140
rect 886 1139 895 1709
rect 855 1130 895 1139
rect 955 1710 995 1720
rect 955 1140 965 1710
rect 985 1140 995 1710
rect 955 1130 995 1140
rect 1055 1710 1095 1720
rect 1055 1140 1065 1710
rect 1085 1140 1095 1710
rect 1055 1130 1095 1140
rect 1155 1710 1195 1720
rect 1155 1140 1165 1710
rect 1185 1140 1195 1710
rect 1155 1130 1195 1140
rect 1255 1710 1295 1720
rect 1255 1140 1265 1710
rect 1285 1140 1295 1710
rect 1255 1130 1295 1140
rect 1355 1710 1395 1720
rect 1355 1140 1365 1710
rect 1385 1140 1395 1710
rect 1355 1130 1395 1140
rect 1455 1710 1495 1720
rect 1455 1140 1465 1710
rect 1485 1140 1495 1710
rect 1455 1130 1495 1140
rect 1555 1710 1595 1720
rect 1555 1139 1565 1710
rect 1585 1139 1595 1710
rect 1555 1130 1595 1139
rect 1614 1709 1645 1720
rect 1614 1137 1620 1709
rect 1640 1137 1645 1709
rect 1614 1130 1645 1137
rect 260 1090 285 1130
rect 460 1090 485 1130
rect 1064 1090 1085 1130
rect 1264 1090 1285 1130
rect 1340 1090 1690 1093
rect 255 1079 1690 1090
rect 255 1072 1350 1079
rect 1341 1055 1350 1072
rect 1370 1074 1690 1079
rect 1370 1055 1380 1074
rect 1341 1045 1380 1055
rect 170 828 209 830
rect -152 820 209 828
rect -152 803 180 820
rect 170 796 180 803
rect 200 803 209 820
rect 200 796 1295 803
rect 170 787 1295 796
rect -195 766 76 786
rect 203 785 1295 787
rect 55 745 75 766
rect 265 745 286 785
rect 465 745 486 785
rect 1065 745 1090 785
rect 1265 745 1290 785
rect -95 737 -64 745
rect -223 635 -178 646
rect -223 616 -215 635
rect -186 619 -178 635
rect -186 616 -149 619
rect -223 608 -149 616
rect -191 50 -149 608
rect -95 166 -90 737
rect -70 166 -64 737
rect -95 155 -64 166
rect -45 735 -5 745
rect -45 165 -35 735
rect -15 165 -5 735
rect -45 155 -5 165
rect 55 735 95 745
rect 55 165 65 735
rect 85 165 95 735
rect 55 155 95 165
rect 155 735 195 745
rect 155 165 165 735
rect 185 165 195 735
rect 155 155 195 165
rect 255 735 295 745
rect 255 165 265 735
rect 285 165 295 735
rect 255 155 295 165
rect 355 735 395 745
rect 355 165 365 735
rect 385 165 395 735
rect 355 155 395 165
rect 455 735 495 745
rect 455 165 465 735
rect 485 165 495 735
rect 455 155 495 165
rect 555 735 595 745
rect 555 165 565 735
rect 585 165 595 735
rect 555 155 595 165
rect 655 735 695 745
rect 655 165 665 735
rect 686 165 695 735
rect 655 155 695 165
rect 755 735 795 745
rect 755 165 765 735
rect 785 165 795 735
rect 755 155 795 165
rect 855 735 895 745
rect 855 734 865 735
rect 855 164 863 734
rect 885 165 895 735
rect 883 164 895 165
rect 855 155 895 164
rect 955 735 995 745
rect 955 165 965 735
rect 985 165 995 735
rect 955 155 995 165
rect 1055 735 1095 745
rect 1055 165 1065 735
rect 1085 165 1095 735
rect 1055 155 1095 165
rect 1155 735 1195 745
rect 1155 165 1165 735
rect 1185 165 1195 735
rect 1155 155 1195 165
rect 1255 735 1295 745
rect 1255 165 1265 735
rect 1285 165 1295 735
rect 1255 155 1295 165
rect 1355 735 1395 745
rect 1355 165 1365 735
rect 1385 165 1395 735
rect 1355 155 1395 165
rect 1455 735 1495 745
rect 1455 165 1465 735
rect 1485 165 1495 735
rect 1455 155 1495 165
rect 1555 735 1595 745
rect 1555 165 1565 735
rect 1585 734 1595 735
rect 1555 164 1566 165
rect 1586 164 1595 734
rect 1555 155 1595 164
rect 1614 735 1645 745
rect 1614 164 1620 735
rect 1640 734 1645 735
rect 1641 164 1645 734
rect 1614 155 1645 164
rect 60 110 80 155
rect 165 151 185 155
rect 100 125 150 135
rect 100 110 110 125
rect 60 100 110 110
rect 140 100 150 125
rect 168 128 185 151
rect 360 128 391 155
rect 565 128 595 155
rect 168 111 595 128
rect 756 110 780 155
rect 956 130 981 155
rect 1155 130 1180 155
rect 1360 130 1383 155
rect 956 110 1383 130
rect 1400 125 1450 135
rect 60 90 150 100
rect 637 91 780 110
rect 637 50 655 91
rect 756 90 780 91
rect 1400 100 1410 125
rect 1440 110 1450 125
rect 1467 110 1487 155
rect 1440 100 1487 110
rect 1400 90 1487 100
rect 1670 70 1689 1074
rect 1736 948 1755 1805
rect 1775 987 1810 995
rect 1775 969 1782 987
rect 1801 969 1810 987
rect 1775 959 1810 969
rect 1706 935 1753 948
rect 1706 915 1724 935
rect 1745 915 1753 935
rect 1706 907 1753 915
rect 1779 829 1796 959
rect -191 31 655 50
rect 637 30 655 31
rect 755 51 1689 70
rect 1773 819 1796 829
rect 1773 818 1793 819
rect -95 -15 -64 -5
rect -95 -587 -90 -15
rect -70 -587 -64 -15
rect -95 -595 -64 -587
rect -45 -15 -5 -5
rect -45 -585 -35 -15
rect -15 -585 -5 -15
rect -45 -595 -5 -585
rect 55 -15 95 -5
rect 55 -585 65 -15
rect 85 -585 95 -15
rect 55 -595 95 -585
rect 155 -15 195 -5
rect 155 -586 165 -15
rect 185 -586 195 -15
rect 155 -595 195 -586
rect 255 -15 295 -5
rect 255 -585 265 -15
rect 285 -585 295 -15
rect 255 -595 295 -585
rect 355 -15 395 -5
rect 355 -585 365 -15
rect 385 -585 395 -15
rect 355 -595 395 -585
rect 455 -15 495 -5
rect 455 -585 465 -15
rect 485 -585 495 -15
rect 455 -595 495 -585
rect 555 -15 595 -5
rect 555 -585 565 -15
rect 585 -585 595 -15
rect 555 -595 595 -585
rect 655 -15 695 -5
rect 655 -585 665 -15
rect 685 -585 695 -15
rect 655 -595 695 -585
rect 755 -15 795 51
rect 755 -585 765 -15
rect 785 -585 795 -15
rect 755 -595 795 -585
rect 855 -15 895 -5
rect 855 -585 865 -15
rect 885 -585 895 -15
rect 855 -595 895 -585
rect 955 -15 995 -5
rect 955 -585 965 -15
rect 985 -585 995 -15
rect 955 -595 995 -585
rect 1055 -15 1095 -5
rect 1055 -585 1065 -15
rect 1085 -585 1095 -15
rect 1055 -595 1095 -585
rect 1155 -15 1195 -5
rect 1155 -585 1165 -15
rect 1185 -585 1195 -15
rect 1155 -595 1195 -585
rect 1255 -15 1295 -5
rect 1255 -585 1265 -15
rect 1285 -585 1295 -15
rect 1255 -595 1295 -585
rect 1355 -15 1395 -5
rect 1355 -588 1365 -15
rect 1385 -588 1395 -15
rect 1355 -595 1395 -588
rect 1455 -15 1495 -5
rect 1455 -585 1465 -15
rect 1485 -585 1495 -15
rect 1455 -595 1495 -585
rect 1555 -15 1595 -5
rect 1555 -585 1565 -15
rect 1585 -585 1595 -15
rect 1555 -595 1595 -585
rect 1614 -14 1645 -5
rect 1614 -585 1620 -14
rect 1640 -585 1645 -14
rect 1614 -595 1645 -585
rect 0 -625 50 -615
rect 0 -645 10 -625
rect 40 -626 50 -625
rect 41 -645 50 -626
rect 0 -654 50 -645
rect 67 -681 93 -595
rect 666 -681 1344 -680
rect 1456 -681 1476 -595
rect 1500 -625 1550 -615
rect 1500 -645 1510 -625
rect 1540 -645 1550 -625
rect 1500 -655 1550 -645
rect 1773 -681 1792 818
rect 65 -699 1792 -681
rect 65 -700 743 -699
rect 1315 -700 1792 -699
<< viali >>
rect 10 2501 40 2520
rect -90 1890 -70 2460
rect 1510 2500 1540 2520
rect -35 1890 -15 2460
rect 165 2460 185 2461
rect 165 1891 185 2460
rect 1366 1890 1385 2459
rect 1385 1890 1386 2459
rect 1366 1889 1386 1890
rect 1565 1890 1585 2460
rect 1620 1890 1640 2460
rect -90 1140 -70 1709
rect -90 1139 -70 1140
rect -35 1140 -15 1710
rect 666 1140 685 1709
rect 685 1140 686 1709
rect 666 1139 686 1140
rect 866 1140 885 1709
rect 885 1140 886 1709
rect 866 1139 886 1140
rect 1565 1140 1585 1709
rect 1565 1139 1585 1140
rect 1620 1138 1640 1707
rect 1620 1137 1640 1138
rect -90 167 -70 737
rect -35 165 -15 735
rect 666 165 685 735
rect 685 165 686 735
rect 863 165 865 734
rect 865 165 883 734
rect 863 164 883 165
rect 1566 165 1585 734
rect 1585 165 1586 734
rect 1566 164 1586 165
rect 1621 164 1640 734
rect 1640 164 1641 734
rect -90 -586 -70 -17
rect -90 -587 -70 -586
rect -35 -585 -15 -15
rect 165 -585 185 -16
rect 165 -586 185 -585
rect 1365 -585 1385 -18
rect 1365 -588 1385 -585
rect 1565 -585 1585 -15
rect 1620 -585 1640 -15
rect 11 -645 40 -626
rect 40 -645 41 -626
rect 1510 -645 1540 -625
<< metal1 >>
rect -198 2520 1765 2537
rect -198 2501 10 2520
rect 40 2501 1510 2520
rect -198 2500 1510 2501
rect 1540 2500 1765 2520
rect -198 2461 1765 2500
rect -198 2460 165 2461
rect -198 1890 -90 2460
rect -70 1890 -35 2460
rect -15 1891 165 2460
rect 185 2460 1765 2461
rect 185 2459 1565 2460
rect 185 1891 1366 2459
rect -15 1890 1366 1891
rect -198 1889 1366 1890
rect 1386 1890 1565 2459
rect 1585 1890 1620 2460
rect 1640 1890 1765 2460
rect 1386 1889 1765 1890
rect -198 1710 1765 1889
rect -198 1709 -35 1710
rect -198 1139 -90 1709
rect -70 1140 -35 1709
rect -15 1709 1765 1710
rect -15 1140 666 1709
rect -70 1139 666 1140
rect 686 1139 866 1709
rect 886 1139 1565 1709
rect 1585 1707 1765 1709
rect 1585 1139 1620 1707
rect -198 1137 1620 1139
rect 1640 1137 1765 1707
rect -198 1038 1765 1137
rect -243 737 1720 848
rect -243 167 -90 737
rect -70 735 1720 737
rect -70 167 -35 735
rect -243 165 -35 167
rect -15 165 666 735
rect 686 734 1720 735
rect 686 165 863 734
rect -243 164 863 165
rect 883 164 1566 734
rect 1586 164 1621 734
rect 1641 164 1720 734
rect -243 -15 1720 164
rect -243 -17 -35 -15
rect -243 -587 -90 -17
rect -70 -585 -35 -17
rect -15 -16 1565 -15
rect -15 -585 165 -16
rect -70 -586 165 -585
rect 185 -18 1565 -16
rect 185 -586 1365 -18
rect -70 -587 1365 -586
rect -243 -588 1365 -587
rect 1385 -585 1565 -18
rect 1585 -585 1620 -15
rect 1640 -585 1720 -15
rect 1385 -588 1720 -585
rect -243 -625 1720 -588
rect -243 -626 1510 -625
rect -243 -645 11 -626
rect 41 -645 1510 -626
rect 1540 -645 1720 -625
rect -243 -661 1720 -645
<< labels >>
rlabel metal1 1763 2521 1763 2521 1 VP
port 2 n
rlabel poly 1818 982 1818 982 1 VCp
port 3 n
rlabel poly 1806 874 1806 874 1 VCn
port 4 n
rlabel metal1 1717 809 1717 809 1 VN
port 6 n
rlabel poly -242 -693 -242 -693 1 VBn
port 5 n
rlabel poly 1999 2611 1999 2611 7 VBp
port 1 w
<< end >>
