magic
tech sky130A
timestamp 1697429884
<< nwell >>
rect 2011 1796 2441 2533
<< poly >>
rect 2248 2576 2307 3339
rect 2248 2550 2386 2576
rect 2342 2549 2386 2550
rect 2298 1794 2376 1818
rect 2298 1699 2324 1794
rect 2093 1680 2324 1699
rect 2081 1678 2324 1680
rect 2078 1575 2143 1594
rect 2107 253 2143 1575
rect 2107 244 2144 253
rect 2108 161 2144 244
rect 2219 238 2269 239
rect 2219 231 2376 238
rect 2219 206 2228 231
rect 2252 216 2376 231
rect 2252 206 2269 216
rect 2219 198 2269 206
rect 2107 120 2366 161
rect 1676 -23 1728 93
rect 1676 -52 1685 -23
rect 1713 -52 1728 -23
rect 1676 -63 1728 -52
<< polycont >>
rect 2228 206 2252 231
rect 1685 -52 1713 -23
<< locali >>
rect 2219 231 2269 240
rect 2219 206 2228 231
rect 2252 206 2269 231
rect 2219 199 2269 206
rect 1676 -22 1728 -11
rect 2220 -22 2269 199
rect 1676 -23 2269 -22
rect 1676 -52 1685 -23
rect 1713 -52 2269 -23
rect 1676 -56 2269 -52
rect 1676 -63 1728 -56
<< metal1 >>
rect 2011 1796 2441 2533
rect 1994 47 2398 1556
use amp  amp_0
timestamp 1697428877
transform 1 0 2455 0 1 84
box -90 -684 1257 2496
use bias  bias_0
timestamp 1697429042
transform 1 0 277 0 1 709
box -277 -709 2001 2630
<< end >>
